magic
tech sky130A
magscale 1 2
timestamp 1671749968
<< viali >>
rect 1685 57545 1719 57579
rect 4077 57545 4111 57579
rect 9873 57545 9907 57579
rect 15669 57545 15703 57579
rect 22109 57545 22143 57579
rect 27261 57545 27295 57579
rect 38301 57545 38335 57579
rect 43361 57545 43395 57579
rect 49157 57545 49191 57579
rect 55689 57545 55723 57579
rect 58265 57545 58299 57579
rect 37565 57477 37599 57511
rect 1869 57409 1903 57443
rect 4261 57409 4295 57443
rect 10057 57409 10091 57443
rect 10517 57409 10551 57443
rect 15853 57409 15887 57443
rect 22293 57409 22327 57443
rect 27445 57409 27479 57443
rect 31769 57409 31803 57443
rect 32321 57409 32355 57443
rect 38117 57409 38151 57443
rect 43545 57409 43579 57443
rect 49341 57409 49375 57443
rect 55505 57409 55539 57443
rect 58081 57409 58115 57443
rect 32505 57341 32539 57375
rect 2329 57205 2363 57239
rect 4721 57205 4755 57239
rect 22753 57205 22787 57239
rect 27997 57205 28031 57239
rect 44005 57205 44039 57239
rect 57529 57205 57563 57239
rect 41153 56797 41187 56831
rect 41797 56797 41831 56831
rect 15945 56661 15979 56695
rect 41337 56661 41371 56695
rect 49433 56661 49467 56695
rect 58081 54621 58115 54655
rect 57529 54485 57563 54519
rect 58265 54485 58299 54519
rect 1869 53533 1903 53567
rect 1685 53397 1719 53431
rect 2421 53397 2455 53431
rect 58081 48705 58115 48739
rect 57529 48501 57563 48535
rect 58265 48501 58299 48535
rect 1685 47141 1719 47175
rect 1869 47005 1903 47039
rect 2421 46937 2455 46971
rect 58081 42653 58115 42687
rect 57529 42517 57563 42551
rect 58265 42517 58299 42551
rect 1869 41089 1903 41123
rect 2329 41089 2363 41123
rect 1685 40885 1719 40919
rect 58081 37213 58115 37247
rect 58265 37077 58299 37111
rect 1869 35649 1903 35683
rect 2329 35649 2363 35683
rect 1685 35445 1719 35479
rect 44833 31297 44867 31331
rect 45201 31297 45235 31331
rect 46765 31297 46799 31331
rect 47041 31297 47075 31331
rect 44281 31093 44315 31127
rect 46949 31093 46983 31127
rect 48421 30753 48455 30787
rect 49249 30753 49283 30787
rect 46305 30685 46339 30719
rect 46949 30685 46983 30719
rect 58081 30685 58115 30719
rect 45753 30617 45787 30651
rect 58265 30549 58299 30583
rect 46213 30345 46247 30379
rect 44833 30277 44867 30311
rect 46121 30277 46155 30311
rect 46581 30277 46615 30311
rect 49801 30277 49835 30311
rect 46397 30209 46431 30243
rect 49617 30209 49651 30243
rect 45293 30141 45327 30175
rect 45109 30073 45143 30107
rect 49433 30005 49467 30039
rect 46765 29801 46799 29835
rect 47317 29801 47351 29835
rect 48789 29801 48823 29835
rect 48145 29733 48179 29767
rect 48973 29733 49007 29767
rect 52009 29733 52043 29767
rect 45661 29665 45695 29699
rect 45845 29665 45879 29699
rect 48329 29665 48363 29699
rect 49249 29665 49283 29699
rect 50905 29665 50939 29699
rect 51549 29665 51583 29699
rect 1869 29597 1903 29631
rect 45569 29597 45603 29631
rect 46305 29597 46339 29631
rect 46581 29597 46615 29631
rect 47225 29597 47259 29631
rect 50813 29597 50847 29631
rect 50997 29597 51031 29631
rect 51641 29597 51675 29631
rect 47869 29529 47903 29563
rect 1685 29461 1719 29495
rect 2421 29461 2455 29495
rect 45201 29461 45235 29495
rect 46397 29461 46431 29495
rect 45293 29257 45327 29291
rect 46137 29257 46171 29291
rect 46305 29257 46339 29291
rect 51825 29257 51859 29291
rect 45937 29189 45971 29223
rect 51641 29189 51675 29223
rect 44649 29121 44683 29155
rect 46765 29121 46799 29155
rect 47961 29121 47995 29155
rect 49249 29121 49283 29155
rect 49709 29121 49743 29155
rect 49985 29121 50019 29155
rect 50353 29121 50387 29155
rect 50721 29121 50755 29155
rect 51457 29121 51491 29155
rect 53849 29121 53883 29155
rect 54493 29121 54527 29155
rect 44741 29053 44775 29087
rect 48421 29053 48455 29087
rect 53021 28985 53055 29019
rect 46121 28917 46155 28951
rect 46857 28917 46891 28951
rect 47225 28917 47259 28951
rect 48145 28917 48179 28951
rect 50997 28917 51031 28951
rect 46213 28713 46247 28747
rect 46765 28713 46799 28747
rect 47225 28713 47259 28747
rect 45983 28645 46017 28679
rect 49801 28645 49835 28679
rect 46121 28577 46155 28611
rect 46857 28577 46891 28611
rect 50721 28577 50755 28611
rect 45845 28509 45879 28543
rect 46305 28509 46339 28543
rect 47041 28509 47075 28543
rect 49249 28509 49283 28543
rect 49433 28509 49467 28543
rect 49617 28509 49651 28543
rect 50537 28509 50571 28543
rect 51365 28509 51399 28543
rect 51549 28509 51583 28543
rect 51917 28509 51951 28543
rect 52285 28509 52319 28543
rect 52929 28509 52963 28543
rect 53665 28509 53699 28543
rect 53849 28509 53883 28543
rect 56793 28509 56827 28543
rect 56977 28509 57011 28543
rect 46765 28441 46799 28475
rect 49525 28441 49559 28475
rect 50353 28373 50387 28407
rect 53021 28373 53055 28407
rect 53849 28373 53883 28407
rect 56977 28373 57011 28407
rect 46581 28169 46615 28203
rect 46305 28101 46339 28135
rect 54769 28101 54803 28135
rect 44649 28033 44683 28067
rect 45109 28033 45143 28067
rect 46213 28033 46247 28067
rect 46397 28033 46431 28067
rect 47869 28033 47903 28067
rect 47961 28033 47995 28067
rect 48513 28033 48547 28067
rect 49341 28033 49375 28067
rect 49709 28033 49743 28067
rect 50353 28033 50387 28067
rect 51181 28033 51215 28067
rect 51365 28033 51399 28067
rect 52193 28033 52227 28067
rect 52377 28033 52411 28067
rect 52929 28033 52963 28067
rect 53297 28033 53331 28067
rect 54033 28033 54067 28067
rect 54401 28033 54435 28067
rect 54677 28033 54711 28067
rect 55873 28033 55907 28067
rect 56149 28033 56183 28067
rect 48329 27965 48363 27999
rect 49801 27965 49835 27999
rect 51089 27965 51123 27999
rect 51273 27965 51307 27999
rect 51549 27965 51583 27999
rect 55229 27965 55263 27999
rect 46029 27897 46063 27931
rect 47133 27829 47167 27863
rect 52285 27829 52319 27863
rect 46121 27625 46155 27659
rect 47225 27625 47259 27659
rect 49249 27625 49283 27659
rect 51089 27625 51123 27659
rect 46857 27557 46891 27591
rect 48237 27557 48271 27591
rect 53757 27557 53791 27591
rect 55597 27557 55631 27591
rect 44649 27489 44683 27523
rect 45937 27489 45971 27523
rect 47777 27489 47811 27523
rect 52285 27489 52319 27523
rect 52929 27489 52963 27523
rect 43913 27421 43947 27455
rect 44005 27421 44039 27455
rect 44189 27421 44223 27455
rect 45753 27421 45787 27455
rect 45845 27421 45879 27455
rect 46121 27421 46155 27455
rect 47041 27421 47075 27455
rect 47225 27421 47259 27455
rect 47869 27421 47903 27455
rect 49433 27421 49467 27455
rect 49709 27421 49743 27455
rect 50629 27421 50663 27455
rect 50905 27421 50939 27455
rect 52377 27421 52411 27455
rect 53665 27421 53699 27455
rect 53849 27421 53883 27455
rect 53941 27421 53975 27455
rect 54125 27421 54159 27455
rect 54585 27421 54619 27455
rect 55505 27421 55539 27455
rect 56977 27421 57011 27455
rect 57897 27421 57931 27455
rect 56425 27353 56459 27387
rect 49617 27285 49651 27319
rect 50721 27285 50755 27319
rect 54677 27285 54711 27319
rect 45937 27081 45971 27115
rect 47777 27081 47811 27115
rect 51181 27081 51215 27115
rect 52377 27081 52411 27115
rect 54401 27081 54435 27115
rect 56057 27081 56091 27115
rect 43545 27013 43579 27047
rect 47961 27013 47995 27047
rect 49801 27013 49835 27047
rect 50813 27013 50847 27047
rect 51013 27013 51047 27047
rect 52929 27013 52963 27047
rect 43453 26945 43487 26979
rect 43729 26945 43763 26979
rect 44189 26945 44223 26979
rect 44833 26945 44867 26979
rect 46213 26945 46247 26979
rect 48053 26945 48087 26979
rect 48145 26945 48179 26979
rect 49709 26945 49743 26979
rect 52193 26945 52227 26979
rect 52377 26945 52411 26979
rect 54309 26945 54343 26979
rect 55229 26945 55263 26979
rect 55413 26945 55447 26979
rect 55873 26945 55907 26979
rect 56057 26945 56091 26979
rect 57069 26945 57103 26979
rect 57161 26945 57195 26979
rect 44925 26877 44959 26911
rect 45937 26877 45971 26911
rect 46673 26877 46707 26911
rect 48329 26877 48363 26911
rect 57253 26877 57287 26911
rect 57345 26877 57379 26911
rect 43729 26809 43763 26843
rect 53205 26809 53239 26843
rect 45477 26741 45511 26775
rect 46121 26741 46155 26775
rect 50997 26741 51031 26775
rect 53389 26741 53423 26775
rect 55229 26741 55263 26775
rect 57529 26741 57563 26775
rect 44097 26537 44131 26571
rect 44281 26537 44315 26571
rect 45661 26537 45695 26571
rect 46305 26537 46339 26571
rect 47041 26537 47075 26571
rect 47777 26537 47811 26571
rect 49617 26537 49651 26571
rect 50905 26537 50939 26571
rect 38853 26469 38887 26503
rect 47317 26469 47351 26503
rect 53021 26469 53055 26503
rect 46397 26401 46431 26435
rect 47041 26401 47075 26435
rect 47961 26401 47995 26435
rect 57897 26401 57931 26435
rect 45385 26333 45419 26367
rect 45477 26333 45511 26367
rect 46489 26333 46523 26367
rect 46949 26333 46983 26367
rect 47777 26333 47811 26367
rect 48145 26333 48179 26367
rect 48789 26333 48823 26367
rect 49157 26333 49191 26367
rect 49249 26333 49283 26367
rect 50629 26333 50663 26367
rect 50721 26333 50755 26367
rect 53849 26333 53883 26367
rect 54033 26333 54067 26367
rect 56241 26333 56275 26367
rect 56517 26333 56551 26367
rect 57989 26333 58023 26367
rect 58265 26333 58299 26367
rect 38485 26265 38519 26299
rect 44265 26265 44299 26299
rect 44465 26265 44499 26299
rect 48053 26265 48087 26299
rect 49617 26265 49651 26299
rect 50905 26265 50939 26299
rect 38945 26197 38979 26231
rect 46121 26197 46155 26231
rect 44649 25993 44683 26027
rect 46121 25993 46155 26027
rect 46857 25993 46891 26027
rect 54033 25993 54067 26027
rect 45201 25925 45235 25959
rect 45753 25925 45787 25959
rect 45958 25925 45992 25959
rect 49157 25925 49191 25959
rect 57253 25925 57287 25959
rect 58173 25925 58207 25959
rect 38945 25857 38979 25891
rect 39037 25857 39071 25891
rect 44005 25857 44039 25891
rect 45293 25857 45327 25891
rect 46581 25857 46615 25891
rect 46673 25857 46707 25891
rect 49433 25857 49467 25891
rect 50353 25857 50387 25891
rect 50721 25857 50755 25891
rect 50997 25857 51031 25891
rect 52929 25857 52963 25891
rect 54033 25857 54067 25891
rect 54217 25857 54251 25891
rect 54953 25857 54987 25891
rect 55045 25857 55079 25891
rect 56057 25857 56091 25891
rect 57069 25857 57103 25891
rect 57161 25857 57195 25891
rect 57437 25857 57471 25891
rect 57529 25857 57563 25891
rect 58081 25857 58115 25891
rect 43913 25789 43947 25823
rect 46857 25789 46891 25823
rect 49249 25789 49283 25823
rect 50813 25789 50847 25823
rect 53021 25789 53055 25823
rect 54769 25789 54803 25823
rect 56149 25789 56183 25823
rect 49617 25721 49651 25755
rect 56425 25721 56459 25755
rect 38117 25653 38151 25687
rect 45937 25653 45971 25687
rect 47777 25653 47811 25687
rect 48329 25653 48363 25687
rect 49157 25653 49191 25687
rect 52929 25653 52963 25687
rect 53297 25653 53331 25687
rect 56057 25653 56091 25687
rect 56885 25653 56919 25687
rect 40417 25449 40451 25483
rect 43913 25449 43947 25483
rect 45477 25449 45511 25483
rect 46213 25449 46247 25483
rect 47501 25449 47535 25483
rect 48789 25449 48823 25483
rect 50813 25449 50847 25483
rect 53941 25449 53975 25483
rect 55965 25449 55999 25483
rect 56057 25449 56091 25483
rect 38945 25381 38979 25415
rect 37269 25313 37303 25347
rect 38393 25313 38427 25347
rect 45385 25313 45419 25347
rect 47317 25313 47351 25347
rect 48605 25313 48639 25347
rect 49341 25313 49375 25347
rect 50629 25313 50663 25347
rect 52193 25313 52227 25347
rect 52837 25313 52871 25347
rect 56149 25313 56183 25347
rect 58081 25313 58115 25347
rect 37473 25245 37507 25279
rect 38025 25245 38059 25279
rect 38209 25245 38243 25279
rect 38853 25245 38887 25279
rect 39221 25245 39255 25279
rect 39405 25245 39439 25279
rect 40049 25245 40083 25279
rect 40233 25245 40267 25279
rect 43729 25245 43763 25279
rect 43913 25245 43947 25279
rect 45753 25245 45787 25279
rect 47225 25245 47259 25279
rect 48513 25245 48547 25279
rect 49525 25245 49559 25279
rect 49801 25245 49835 25279
rect 50537 25245 50571 25279
rect 52929 25245 52963 25279
rect 53941 25245 53975 25279
rect 54125 25245 54159 25279
rect 55873 25245 55907 25279
rect 37197 25177 37231 25211
rect 57253 25177 57287 25211
rect 37381 25109 37415 25143
rect 44373 25109 44407 25143
rect 45569 25109 45603 25143
rect 45661 25109 45695 25143
rect 49709 25109 49743 25143
rect 56793 25109 56827 25143
rect 36461 24905 36495 24939
rect 37673 24905 37707 24939
rect 37841 24905 37875 24939
rect 38761 24905 38795 24939
rect 40233 24905 40267 24939
rect 47777 24905 47811 24939
rect 48989 24905 49023 24939
rect 50537 24905 50571 24939
rect 37473 24837 37507 24871
rect 44649 24837 44683 24871
rect 46397 24837 46431 24871
rect 48789 24837 48823 24871
rect 35173 24769 35207 24803
rect 36093 24769 36127 24803
rect 38669 24769 38703 24803
rect 38945 24769 38979 24803
rect 40141 24769 40175 24803
rect 40325 24769 40359 24803
rect 43821 24769 43855 24803
rect 45661 24769 45695 24803
rect 45753 24769 45787 24803
rect 46673 24769 46707 24803
rect 47961 24769 47995 24803
rect 48145 24769 48179 24803
rect 49709 24769 49743 24803
rect 50169 24769 50203 24803
rect 50261 24769 50295 24803
rect 52193 24769 52227 24803
rect 52377 24769 52411 24803
rect 52929 24769 52963 24803
rect 53021 24769 53055 24803
rect 53205 24769 53239 24803
rect 53389 24769 53423 24803
rect 54769 24769 54803 24803
rect 55505 24769 55539 24803
rect 57069 24769 57103 24803
rect 57253 24769 57287 24803
rect 58081 24769 58115 24803
rect 34897 24701 34931 24735
rect 36185 24701 36219 24735
rect 45569 24701 45603 24735
rect 45845 24701 45879 24735
rect 46397 24701 46431 24735
rect 47133 24701 47167 24735
rect 52285 24701 52319 24735
rect 56425 24701 56459 24735
rect 34989 24633 35023 24667
rect 38945 24633 38979 24667
rect 44281 24633 44315 24667
rect 44833 24633 44867 24667
rect 49157 24633 49191 24667
rect 35357 24565 35391 24599
rect 37657 24565 37691 24599
rect 43821 24565 43855 24599
rect 44649 24565 44683 24599
rect 45385 24565 45419 24599
rect 46581 24565 46615 24599
rect 48973 24565 49007 24599
rect 50169 24565 50203 24599
rect 57161 24565 57195 24599
rect 58265 24565 58299 24599
rect 35449 24361 35483 24395
rect 36737 24361 36771 24395
rect 37105 24361 37139 24395
rect 38393 24361 38427 24395
rect 40049 24361 40083 24395
rect 44005 24361 44039 24395
rect 45385 24361 45419 24395
rect 47593 24361 47627 24395
rect 50537 24361 50571 24395
rect 55873 24361 55907 24395
rect 57161 24361 57195 24395
rect 35357 24225 35391 24259
rect 43269 24225 43303 24259
rect 50905 24225 50939 24259
rect 54953 24225 54987 24259
rect 56793 24225 56827 24259
rect 57621 24225 57655 24259
rect 27537 24157 27571 24191
rect 27721 24157 27755 24191
rect 31953 24157 31987 24191
rect 32505 24157 32539 24191
rect 35265 24157 35299 24191
rect 36645 24157 36679 24191
rect 38393 24157 38427 24191
rect 38577 24157 38611 24191
rect 40233 24157 40267 24191
rect 40601 24157 40635 24191
rect 40693 24157 40727 24191
rect 43177 24157 43211 24191
rect 43361 24157 43395 24191
rect 43821 24157 43855 24191
rect 46581 24157 46615 24191
rect 46857 24157 46891 24191
rect 50813 24157 50847 24191
rect 52653 24157 52687 24191
rect 53849 24157 53883 24191
rect 54217 24157 54251 24191
rect 54677 24157 54711 24191
rect 55505 24157 55539 24191
rect 55689 24157 55723 24191
rect 56701 24157 56735 24191
rect 56977 24157 57011 24191
rect 57805 24157 57839 24191
rect 58081 24157 58115 24191
rect 40325 24089 40359 24123
rect 40417 24089 40451 24123
rect 45369 24089 45403 24123
rect 45569 24089 45603 24123
rect 46765 24089 46799 24123
rect 52469 24089 52503 24123
rect 57989 24089 58023 24123
rect 27629 24021 27663 24055
rect 35633 24021 35667 24055
rect 45201 24021 45235 24055
rect 46857 24021 46891 24055
rect 52837 24021 52871 24055
rect 28825 23817 28859 23851
rect 31585 23817 31619 23851
rect 34989 23817 35023 23851
rect 36369 23817 36403 23851
rect 38761 23817 38795 23851
rect 39957 23817 39991 23851
rect 44649 23817 44683 23851
rect 45937 23817 45971 23851
rect 47977 23817 48011 23851
rect 48145 23817 48179 23851
rect 49893 23817 49927 23851
rect 50813 23817 50847 23851
rect 53113 23817 53147 23851
rect 54217 23817 54251 23851
rect 56425 23817 56459 23851
rect 58173 23817 58207 23851
rect 38945 23749 38979 23783
rect 47777 23749 47811 23783
rect 48605 23749 48639 23783
rect 48821 23749 48855 23783
rect 50445 23749 50479 23783
rect 52377 23749 52411 23783
rect 1869 23681 1903 23715
rect 2329 23681 2363 23715
rect 25605 23681 25639 23715
rect 27813 23681 27847 23715
rect 27997 23681 28031 23715
rect 30205 23681 30239 23715
rect 31401 23681 31435 23715
rect 31585 23681 31619 23715
rect 35265 23681 35299 23715
rect 35909 23681 35943 23715
rect 36369 23681 36403 23715
rect 36553 23681 36587 23715
rect 39129 23681 39163 23715
rect 40234 23681 40268 23715
rect 40417 23681 40451 23715
rect 40969 23681 41003 23715
rect 41153 23681 41187 23715
rect 42625 23681 42659 23715
rect 42809 23681 42843 23715
rect 43913 23681 43947 23715
rect 44465 23681 44499 23715
rect 45201 23681 45235 23715
rect 45385 23681 45419 23715
rect 46673 23681 46707 23715
rect 46765 23681 46799 23715
rect 46949 23681 46983 23715
rect 49709 23681 49743 23715
rect 50629 23681 50663 23715
rect 51273 23681 51307 23715
rect 51457 23681 51491 23715
rect 52101 23681 52135 23715
rect 52193 23681 52227 23715
rect 53021 23681 53055 23715
rect 53205 23681 53239 23715
rect 53849 23681 53883 23715
rect 56333 23681 56367 23715
rect 56517 23681 56551 23715
rect 58357 23681 58391 23715
rect 24593 23613 24627 23647
rect 30021 23613 30055 23647
rect 34989 23613 35023 23647
rect 40141 23613 40175 23647
rect 40325 23613 40359 23647
rect 45293 23613 45327 23647
rect 49433 23613 49467 23647
rect 53941 23613 53975 23647
rect 57069 23613 57103 23647
rect 30389 23545 30423 23579
rect 57345 23545 57379 23579
rect 1685 23477 1719 23511
rect 35173 23477 35207 23511
rect 35817 23477 35851 23511
rect 41061 23477 41095 23511
rect 41705 23477 41739 23511
rect 42717 23477 42751 23511
rect 43821 23477 43855 23511
rect 47133 23477 47167 23511
rect 47961 23477 47995 23511
rect 48789 23477 48823 23511
rect 48973 23477 49007 23511
rect 49525 23477 49559 23511
rect 51641 23477 51675 23511
rect 52377 23477 52411 23511
rect 57529 23477 57563 23511
rect 28457 23273 28491 23307
rect 29745 23273 29779 23307
rect 34253 23273 34287 23307
rect 35357 23273 35391 23307
rect 38577 23273 38611 23307
rect 39037 23273 39071 23307
rect 43453 23273 43487 23307
rect 45661 23273 45695 23307
rect 46489 23273 46523 23307
rect 48973 23273 49007 23307
rect 49801 23273 49835 23307
rect 52101 23273 52135 23307
rect 52285 23273 52319 23307
rect 53573 23273 53607 23307
rect 53757 23273 53791 23307
rect 57621 23273 57655 23307
rect 58265 23273 58299 23307
rect 28641 23205 28675 23239
rect 44649 23205 44683 23239
rect 45293 23205 45327 23239
rect 49709 23205 49743 23239
rect 50353 23205 50387 23239
rect 56057 23205 56091 23239
rect 26157 23137 26191 23171
rect 31125 23137 31159 23171
rect 36369 23137 36403 23171
rect 36645 23137 36679 23171
rect 37381 23137 37415 23171
rect 37657 23137 37691 23171
rect 41981 23137 42015 23171
rect 44373 23137 44407 23171
rect 47685 23137 47719 23171
rect 48145 23137 48179 23171
rect 55597 23137 55631 23171
rect 23121 23069 23155 23103
rect 23581 23069 23615 23103
rect 26065 23069 26099 23103
rect 26709 23069 26743 23103
rect 27077 23069 27111 23103
rect 27445 23069 27479 23103
rect 27997 23069 28031 23103
rect 29929 23069 29963 23103
rect 30205 23069 30239 23103
rect 30757 23069 30791 23103
rect 31033 23069 31067 23103
rect 31677 23069 31711 23103
rect 31769 23069 31803 23103
rect 31861 23069 31895 23103
rect 31953 23069 31987 23103
rect 34161 23069 34195 23103
rect 34345 23069 34379 23103
rect 35173 23069 35207 23103
rect 36277 23069 36311 23103
rect 37289 23069 37323 23103
rect 38117 23069 38151 23103
rect 38209 23069 38243 23103
rect 38393 23069 38427 23103
rect 39037 23069 39071 23103
rect 39129 23069 39163 23103
rect 40509 23069 40543 23103
rect 40877 23069 40911 23103
rect 41705 23069 41739 23103
rect 44281 23069 44315 23103
rect 45569 23069 45603 23103
rect 45661 23069 45695 23103
rect 46305 23069 46339 23103
rect 47777 23069 47811 23103
rect 48697 23069 48731 23103
rect 48973 23069 49007 23103
rect 49801 23069 49835 23103
rect 55689 23069 55723 23103
rect 58081 23069 58115 23103
rect 58265 23069 58299 23103
rect 28917 23001 28951 23035
rect 34989 23001 35023 23035
rect 39313 23001 39347 23035
rect 46121 23001 46155 23035
rect 49525 23001 49559 23035
rect 51917 23001 51951 23035
rect 53389 23001 53423 23035
rect 53605 23001 53639 23035
rect 57253 23001 57287 23035
rect 57437 23001 57471 23035
rect 22753 22933 22787 22967
rect 30113 22933 30147 22967
rect 32137 22933 32171 22967
rect 41245 22933 41279 22967
rect 48789 22933 48823 22967
rect 52117 22933 52151 22967
rect 26617 22729 26651 22763
rect 29009 22729 29043 22763
rect 37841 22729 37875 22763
rect 39405 22729 39439 22763
rect 40509 22729 40543 22763
rect 41981 22729 42015 22763
rect 44373 22729 44407 22763
rect 45937 22729 45971 22763
rect 46581 22729 46615 22763
rect 47961 22729 47995 22763
rect 48053 22729 48087 22763
rect 50997 22729 51031 22763
rect 56977 22729 57011 22763
rect 58173 22729 58207 22763
rect 37657 22661 37691 22695
rect 39313 22661 39347 22695
rect 42901 22661 42935 22695
rect 45477 22661 45511 22695
rect 48145 22661 48179 22695
rect 56609 22661 56643 22695
rect 56809 22661 56843 22695
rect 25973 22593 26007 22627
rect 28825 22593 28859 22627
rect 29469 22593 29503 22627
rect 29929 22593 29963 22627
rect 30297 22593 30331 22627
rect 30665 22593 30699 22627
rect 31033 22593 31067 22627
rect 31309 22593 31343 22627
rect 33977 22593 34011 22627
rect 34805 22593 34839 22627
rect 37473 22593 37507 22627
rect 39129 22593 39163 22627
rect 39405 22593 39439 22627
rect 39865 22593 39899 22627
rect 40509 22593 40543 22627
rect 40693 22593 40727 22627
rect 41153 22593 41187 22627
rect 41337 22593 41371 22627
rect 45753 22593 45787 22627
rect 47777 22593 47811 22627
rect 49341 22593 49375 22627
rect 49525 22593 49559 22627
rect 50629 22593 50663 22627
rect 51733 22593 51767 22627
rect 53389 22593 53423 22627
rect 53573 22593 53607 22627
rect 53849 22593 53883 22627
rect 54125 22593 54159 22627
rect 54217 22593 54251 22627
rect 54953 22593 54987 22627
rect 55137 22593 55171 22627
rect 55597 22593 55631 22627
rect 23581 22525 23615 22559
rect 26065 22525 26099 22559
rect 28549 22525 28583 22559
rect 39957 22525 39991 22559
rect 42625 22525 42659 22559
rect 45661 22525 45695 22559
rect 46029 22525 46063 22559
rect 46121 22525 46155 22559
rect 50537 22525 50571 22559
rect 51641 22525 51675 22559
rect 52101 22525 52135 22559
rect 23305 22457 23339 22491
rect 28641 22457 28675 22491
rect 44925 22457 44959 22491
rect 48329 22457 48363 22491
rect 23121 22389 23155 22423
rect 24961 22389 24995 22423
rect 41245 22389 41279 22423
rect 47225 22389 47259 22423
rect 49525 22389 49559 22423
rect 55045 22389 55079 22423
rect 55689 22389 55723 22423
rect 56057 22389 56091 22423
rect 56793 22389 56827 22423
rect 27537 22185 27571 22219
rect 27997 22185 28031 22219
rect 28365 22185 28399 22219
rect 30757 22185 30791 22219
rect 34897 22185 34931 22219
rect 42717 22185 42751 22219
rect 44465 22185 44499 22219
rect 48881 22185 48915 22219
rect 50813 22185 50847 22219
rect 53297 22185 53331 22219
rect 56793 22185 56827 22219
rect 58173 22185 58207 22219
rect 33333 22117 33367 22151
rect 43637 22117 43671 22151
rect 46765 22117 46799 22151
rect 25053 22049 25087 22083
rect 33793 22049 33827 22083
rect 39497 22049 39531 22083
rect 41981 22049 42015 22083
rect 47225 22049 47259 22083
rect 49249 22049 49283 22083
rect 49341 22049 49375 22083
rect 50445 22049 50479 22083
rect 53573 22049 53607 22083
rect 54401 22049 54435 22083
rect 55873 22049 55907 22083
rect 57805 22049 57839 22083
rect 23949 21981 23983 22015
rect 24041 21981 24075 22015
rect 24869 21981 24903 22015
rect 25973 21981 26007 22015
rect 26341 21981 26375 22015
rect 27077 21981 27111 22015
rect 27169 21981 27203 22015
rect 27353 21981 27387 22015
rect 27997 21981 28031 22015
rect 28089 21981 28123 22015
rect 30941 21981 30975 22015
rect 31125 21981 31159 22015
rect 31217 21981 31251 22015
rect 31677 21981 31711 22015
rect 31769 21981 31803 22015
rect 32045 21981 32079 22015
rect 32137 21981 32171 22015
rect 33701 21981 33735 22015
rect 35541 21981 35575 22015
rect 36369 21981 36403 22015
rect 39037 21981 39071 22015
rect 39313 21981 39347 22015
rect 40693 21981 40727 22015
rect 41061 21981 41095 22015
rect 41153 21981 41187 22015
rect 41705 21981 41739 22015
rect 41797 21981 41831 22015
rect 41889 21981 41923 22015
rect 44189 21981 44223 22015
rect 45845 21981 45879 22015
rect 47133 21981 47167 22015
rect 49065 21981 49099 22015
rect 49157 21981 49191 22015
rect 50537 21981 50571 22015
rect 52469 21981 52503 22015
rect 53481 21981 53515 22015
rect 53665 21981 53699 22015
rect 53757 21981 53791 22015
rect 54309 21981 54343 22015
rect 54493 21981 54527 22015
rect 55689 21981 55723 22015
rect 56517 21981 56551 22015
rect 57897 21981 57931 22015
rect 23765 21913 23799 21947
rect 24593 21913 24627 21947
rect 31953 21913 31987 21947
rect 40785 21913 40819 21947
rect 40877 21913 40911 21947
rect 44465 21913 44499 21947
rect 52653 21913 52687 21947
rect 52837 21913 52871 21947
rect 55505 21913 55539 21947
rect 56793 21913 56827 21947
rect 23863 21845 23897 21879
rect 24685 21845 24719 21879
rect 25973 21845 26007 21879
rect 26157 21845 26191 21879
rect 26249 21845 26283 21879
rect 32321 21845 32355 21879
rect 39129 21845 39163 21879
rect 40509 21845 40543 21879
rect 42165 21845 42199 21879
rect 44281 21845 44315 21879
rect 46029 21845 46063 21879
rect 56609 21845 56643 21879
rect 24501 21641 24535 21675
rect 24869 21641 24903 21675
rect 26341 21641 26375 21675
rect 26617 21641 26651 21675
rect 27721 21641 27755 21675
rect 31769 21641 31803 21675
rect 32597 21641 32631 21675
rect 36645 21641 36679 21675
rect 39037 21641 39071 21675
rect 40601 21641 40635 21675
rect 41245 21641 41279 21675
rect 47777 21641 47811 21675
rect 48789 21641 48823 21675
rect 55137 21641 55171 21675
rect 56977 21641 57011 21675
rect 58173 21641 58207 21675
rect 30573 21573 30607 21607
rect 35725 21573 35759 21607
rect 43729 21573 43763 21607
rect 44833 21573 44867 21607
rect 23305 21505 23339 21539
rect 24685 21505 24719 21539
rect 24961 21505 24995 21539
rect 25605 21505 25639 21539
rect 26249 21505 26283 21539
rect 26433 21505 26467 21539
rect 28089 21505 28123 21539
rect 30021 21505 30055 21539
rect 30481 21505 30515 21539
rect 30665 21505 30699 21539
rect 31677 21505 31711 21539
rect 31769 21505 31803 21539
rect 32321 21505 32355 21539
rect 33701 21505 33735 21539
rect 33885 21505 33919 21539
rect 35357 21505 35391 21539
rect 35541 21505 35575 21539
rect 36461 21505 36495 21539
rect 36645 21505 36679 21539
rect 37657 21505 37691 21539
rect 38669 21505 38703 21539
rect 40509 21505 40543 21539
rect 41153 21505 41187 21539
rect 42717 21505 42751 21539
rect 47777 21505 47811 21539
rect 47961 21505 47995 21539
rect 48973 21505 49007 21539
rect 49341 21505 49375 21539
rect 54125 21505 54159 21539
rect 54401 21505 54435 21539
rect 54585 21505 54619 21539
rect 55045 21505 55079 21539
rect 55229 21505 55263 21539
rect 56885 21505 56919 21539
rect 57069 21505 57103 21539
rect 58081 21505 58115 21539
rect 58265 21505 58299 21539
rect 22477 21437 22511 21471
rect 23397 21437 23431 21471
rect 27997 21437 28031 21471
rect 31493 21437 31527 21471
rect 32597 21437 32631 21471
rect 33149 21437 33183 21471
rect 34437 21437 34471 21471
rect 37565 21437 37599 21471
rect 38025 21437 38059 21471
rect 38577 21437 38611 21471
rect 44557 21437 44591 21471
rect 26065 21369 26099 21403
rect 32413 21369 32447 21403
rect 25513 21301 25547 21335
rect 27261 21301 27295 21335
rect 33793 21301 33827 21335
rect 46305 21301 46339 21335
rect 46949 21301 46983 21335
rect 48973 21301 49007 21335
rect 54217 21301 54251 21335
rect 23673 21097 23707 21131
rect 24593 21097 24627 21131
rect 24777 21097 24811 21131
rect 25973 21097 26007 21131
rect 27813 21097 27847 21131
rect 27997 21097 28031 21131
rect 29837 21097 29871 21131
rect 31493 21097 31527 21131
rect 32321 21097 32355 21131
rect 33149 21097 33183 21131
rect 33333 21097 33367 21131
rect 35909 21097 35943 21131
rect 37565 21097 37599 21131
rect 38577 21097 38611 21131
rect 44649 21097 44683 21131
rect 45845 21097 45879 21131
rect 48881 21097 48915 21131
rect 54125 21097 54159 21131
rect 56885 21097 56919 21131
rect 57713 21097 57747 21131
rect 57897 21097 57931 21131
rect 31677 21029 31711 21063
rect 34161 21029 34195 21063
rect 41521 21029 41555 21063
rect 42349 21029 42383 21063
rect 47501 21029 47535 21063
rect 52561 21029 52595 21063
rect 26249 20961 26283 20995
rect 28549 20961 28583 20995
rect 28733 20961 28767 20995
rect 33977 20961 34011 20995
rect 35633 20961 35667 20995
rect 38209 20961 38243 20995
rect 41981 20961 42015 20995
rect 42901 20961 42935 20995
rect 47225 20961 47259 20995
rect 48053 20961 48087 20995
rect 52101 20961 52135 20995
rect 55597 20961 55631 20995
rect 23857 20893 23891 20927
rect 24041 20893 24075 20927
rect 26157 20893 26191 20927
rect 26341 20893 26375 20927
rect 26433 20893 26467 20927
rect 28457 20893 28491 20927
rect 30021 20893 30055 20927
rect 30205 20893 30239 20927
rect 30297 20893 30331 20927
rect 31401 20893 31435 20927
rect 31493 20893 31527 20927
rect 32229 20893 32263 20927
rect 34161 20893 34195 20927
rect 35541 20893 35575 20927
rect 37381 20893 37415 20927
rect 37565 20893 37599 20927
rect 38393 20893 38427 20927
rect 47133 20893 47167 20927
rect 47961 20893 47995 20927
rect 48145 20893 48179 20927
rect 48697 20893 48731 20927
rect 48881 20893 48915 20927
rect 49157 20893 49191 20927
rect 50997 20893 51031 20927
rect 51365 20893 51399 20927
rect 51549 20893 51583 20927
rect 52193 20893 52227 20927
rect 53021 20893 53055 20927
rect 53113 20893 53147 20927
rect 53297 20893 53331 20927
rect 53941 20893 53975 20927
rect 54309 20893 54343 20927
rect 54401 20893 54435 20927
rect 55735 20893 55769 20927
rect 24761 20825 24795 20859
rect 24961 20825 24995 20859
rect 27629 20825 27663 20859
rect 28733 20825 28767 20859
rect 31217 20825 31251 20859
rect 32965 20825 32999 20859
rect 33181 20825 33215 20859
rect 33793 20825 33827 20859
rect 43177 20825 43211 20859
rect 53481 20825 53515 20859
rect 56517 20825 56551 20859
rect 56701 20825 56735 20859
rect 57529 20825 57563 20859
rect 27829 20757 27863 20791
rect 36461 20757 36495 20791
rect 42441 20757 42475 20791
rect 45201 20757 45235 20791
rect 46305 20757 46339 20791
rect 51089 20757 51123 20791
rect 56057 20757 56091 20791
rect 57729 20757 57763 20791
rect 24317 20553 24351 20587
rect 25697 20553 25731 20587
rect 26249 20553 26283 20587
rect 26433 20553 26467 20587
rect 28089 20553 28123 20587
rect 29101 20553 29135 20587
rect 30481 20553 30515 20587
rect 31493 20553 31527 20587
rect 32505 20553 32539 20587
rect 33793 20553 33827 20587
rect 35081 20553 35115 20587
rect 39221 20553 39255 20587
rect 41061 20553 41095 20587
rect 43361 20553 43395 20587
rect 48421 20553 48455 20587
rect 53205 20553 53239 20587
rect 56057 20553 56091 20587
rect 58173 20553 58207 20587
rect 22845 20485 22879 20519
rect 28641 20485 28675 20519
rect 32689 20485 32723 20519
rect 46765 20485 46799 20519
rect 49341 20485 49375 20519
rect 50353 20485 50387 20519
rect 51641 20485 51675 20519
rect 54769 20485 54803 20519
rect 56701 20485 56735 20519
rect 58357 20485 58391 20519
rect 23581 20417 23615 20451
rect 24593 20417 24627 20451
rect 24685 20417 24719 20451
rect 25513 20417 25547 20451
rect 26525 20417 26559 20451
rect 26617 20417 26651 20451
rect 27905 20417 27939 20451
rect 28089 20417 28123 20451
rect 29469 20417 29503 20451
rect 30481 20417 30515 20451
rect 30665 20417 30699 20451
rect 30941 20417 30975 20451
rect 31401 20417 31435 20451
rect 31677 20417 31711 20451
rect 31769 20417 31803 20451
rect 32597 20417 32631 20451
rect 33333 20417 33367 20451
rect 33425 20417 33459 20451
rect 33609 20417 33643 20451
rect 35449 20417 35483 20451
rect 36645 20417 36679 20451
rect 36829 20417 36863 20451
rect 38853 20417 38887 20451
rect 40233 20417 40267 20451
rect 41521 20417 41555 20451
rect 41705 20417 41739 20451
rect 42625 20417 42659 20451
rect 44465 20417 44499 20451
rect 45845 20417 45879 20451
rect 46029 20417 46063 20451
rect 46581 20417 46615 20451
rect 48237 20417 48271 20451
rect 48881 20417 48915 20451
rect 48973 20417 49007 20451
rect 49249 20417 49283 20451
rect 50077 20417 50111 20451
rect 50169 20417 50203 20451
rect 50997 20417 51031 20451
rect 51181 20417 51215 20451
rect 51457 20417 51491 20451
rect 52929 20417 52963 20451
rect 54125 20417 54159 20451
rect 54309 20417 54343 20451
rect 54401 20417 54435 20451
rect 54510 20417 54544 20451
rect 55597 20417 55631 20451
rect 56609 20417 56643 20451
rect 56793 20417 56827 20451
rect 58081 20417 58115 20451
rect 24501 20349 24535 20383
rect 24777 20349 24811 20383
rect 26249 20349 26283 20383
rect 29377 20349 29411 20383
rect 30803 20349 30837 20383
rect 31585 20349 31619 20383
rect 32321 20349 32355 20383
rect 32873 20349 32907 20383
rect 35541 20349 35575 20383
rect 38761 20349 38795 20383
rect 40325 20349 40359 20383
rect 44373 20349 44407 20383
rect 45661 20349 45695 20383
rect 48053 20349 48087 20383
rect 50353 20349 50387 20383
rect 53205 20349 53239 20383
rect 44833 20281 44867 20315
rect 58357 20281 58391 20315
rect 36093 20213 36127 20247
rect 36829 20213 36863 20247
rect 41705 20213 41739 20247
rect 42809 20213 42843 20247
rect 49157 20213 49191 20247
rect 52101 20213 52135 20247
rect 53021 20213 53055 20247
rect 55689 20213 55723 20247
rect 57253 20213 57287 20247
rect 23489 20009 23523 20043
rect 23949 20009 23983 20043
rect 27077 20009 27111 20043
rect 29745 20009 29779 20043
rect 31585 20009 31619 20043
rect 33517 20009 33551 20043
rect 35265 20009 35299 20043
rect 38117 20009 38151 20043
rect 38853 20009 38887 20043
rect 39221 20009 39255 20043
rect 40417 20009 40451 20043
rect 44373 20009 44407 20043
rect 46949 20009 46983 20043
rect 47409 20009 47443 20043
rect 49157 20009 49191 20043
rect 51641 20009 51675 20043
rect 54493 20009 54527 20043
rect 55781 20009 55815 20043
rect 57805 20009 57839 20043
rect 26525 19941 26559 19975
rect 37197 19941 37231 19975
rect 46581 19941 46615 19975
rect 47685 19941 47719 19975
rect 47777 19941 47811 19975
rect 50905 19941 50939 19975
rect 24593 19873 24627 19907
rect 25513 19873 25547 19907
rect 28273 19873 28307 19907
rect 28457 19873 28491 19907
rect 36553 19873 36587 19907
rect 36737 19873 36771 19907
rect 37933 19873 37967 19907
rect 40049 19873 40083 19907
rect 41429 19873 41463 19907
rect 42809 19873 42843 19907
rect 46489 19873 46523 19907
rect 49157 19873 49191 19907
rect 52285 19873 52319 19907
rect 53297 19873 53331 19907
rect 54401 19873 54435 19907
rect 56609 19873 56643 19907
rect 57437 19873 57471 19907
rect 23765 19805 23799 19839
rect 24041 19805 24075 19839
rect 25329 19805 25363 19839
rect 26801 19805 26835 19839
rect 28365 19805 28399 19839
rect 28542 19805 28576 19839
rect 29929 19805 29963 19839
rect 30021 19805 30055 19839
rect 31493 19805 31527 19839
rect 31677 19805 31711 19839
rect 33333 19805 33367 19839
rect 35633 19805 35667 19839
rect 37841 19805 37875 19839
rect 38761 19805 38795 19839
rect 40233 19805 40267 19839
rect 43085 19805 43119 19839
rect 44281 19805 44315 19839
rect 44465 19805 44499 19839
rect 45569 19805 45603 19839
rect 45753 19805 45787 19839
rect 46765 19805 46799 19839
rect 47593 19805 47627 19839
rect 47869 19805 47903 19839
rect 48881 19805 48915 19839
rect 49065 19805 49099 19839
rect 50445 19805 50479 19839
rect 50997 19805 51031 19839
rect 51089 19805 51123 19839
rect 52009 19805 52043 19839
rect 53021 19805 53055 19839
rect 53205 19805 53239 19839
rect 53389 19805 53423 19839
rect 53481 19805 53515 19839
rect 54125 19805 54159 19839
rect 54217 19805 54251 19839
rect 54493 19805 54527 19839
rect 55505 19805 55539 19839
rect 56425 19805 56459 19839
rect 56701 19805 56735 19839
rect 57529 19805 57563 19839
rect 26893 19737 26927 19771
rect 33425 19737 33459 19771
rect 33609 19737 33643 19771
rect 35449 19737 35483 19771
rect 42257 19737 42291 19771
rect 45937 19737 45971 19771
rect 48789 19737 48823 19771
rect 53665 19737 53699 19771
rect 55781 19737 55815 19771
rect 56241 19737 56275 19771
rect 26709 19669 26743 19703
rect 28089 19669 28123 19703
rect 29101 19669 29135 19703
rect 36829 19669 36863 19703
rect 43821 19669 43855 19703
rect 52101 19669 52135 19703
rect 55597 19669 55631 19703
rect 23765 19465 23799 19499
rect 24685 19465 24719 19499
rect 25513 19465 25547 19499
rect 26065 19465 26099 19499
rect 34897 19465 34931 19499
rect 36921 19465 36955 19499
rect 37933 19465 37967 19499
rect 41245 19465 41279 19499
rect 41889 19465 41923 19499
rect 42809 19465 42843 19499
rect 43729 19465 43763 19499
rect 48145 19465 48179 19499
rect 50629 19465 50663 19499
rect 51365 19465 51399 19499
rect 51733 19465 51767 19499
rect 53113 19465 53147 19499
rect 55119 19465 55153 19499
rect 57161 19465 57195 19499
rect 28825 19397 28859 19431
rect 29561 19397 29595 19431
rect 33609 19397 33643 19431
rect 36461 19397 36495 19431
rect 39405 19397 39439 19431
rect 39865 19397 39899 19431
rect 40065 19397 40099 19431
rect 46673 19397 46707 19431
rect 51825 19397 51859 19431
rect 55597 19397 55631 19431
rect 24409 19329 24443 19363
rect 24777 19329 24811 19363
rect 25421 19329 25455 19363
rect 25605 19329 25639 19363
rect 26433 19329 26467 19363
rect 28089 19329 28123 19363
rect 28733 19329 28767 19363
rect 28917 19329 28951 19363
rect 29929 19329 29963 19363
rect 30021 19329 30055 19363
rect 31585 19329 31619 19363
rect 31769 19329 31803 19363
rect 32597 19329 32631 19363
rect 33425 19329 33459 19363
rect 34253 19329 34287 19363
rect 34437 19329 34471 19363
rect 34713 19335 34747 19369
rect 35357 19329 35391 19363
rect 35541 19329 35575 19363
rect 35817 19329 35851 19363
rect 36001 19329 36035 19363
rect 37841 19329 37875 19363
rect 38025 19329 38059 19363
rect 41153 19329 41187 19363
rect 41797 19329 41831 19363
rect 41981 19329 42015 19363
rect 42625 19329 42659 19363
rect 43637 19329 43671 19363
rect 46029 19329 46063 19363
rect 48237 19329 48271 19363
rect 48789 19329 48823 19363
rect 49065 19329 49099 19363
rect 49341 19329 49375 19363
rect 50169 19329 50203 19363
rect 50261 19329 50295 19363
rect 53389 19329 53423 19363
rect 56793 19329 56827 19363
rect 22017 19261 22051 19295
rect 22293 19261 22327 19295
rect 26249 19261 26283 19295
rect 26341 19261 26375 19295
rect 26525 19261 26559 19295
rect 27721 19261 27755 19295
rect 28181 19261 28215 19295
rect 29745 19261 29779 19295
rect 29837 19261 29871 19295
rect 32505 19261 32539 19295
rect 32965 19261 32999 19295
rect 33793 19261 33827 19295
rect 43913 19261 43947 19295
rect 44465 19261 44499 19295
rect 45017 19261 45051 19295
rect 46121 19261 46155 19295
rect 48969 19261 49003 19295
rect 49985 19261 50019 19295
rect 52009 19261 52043 19295
rect 53113 19261 53147 19295
rect 55505 19261 55539 19295
rect 55689 19261 55723 19295
rect 56701 19261 56735 19295
rect 31401 19193 31435 19227
rect 36737 19193 36771 19227
rect 48881 19193 48915 19227
rect 27169 19125 27203 19159
rect 40049 19125 40083 19159
rect 40233 19125 40267 19159
rect 43269 19125 43303 19159
rect 45753 19125 45787 19159
rect 53297 19125 53331 19159
rect 53849 19125 53883 19159
rect 54401 19125 54435 19159
rect 58173 19125 58207 19159
rect 22109 18921 22143 18955
rect 23857 18921 23891 18955
rect 29101 18921 29135 18955
rect 30757 18921 30791 18955
rect 31585 18921 31619 18955
rect 32505 18921 32539 18955
rect 34897 18921 34931 18955
rect 35173 18921 35207 18955
rect 38209 18921 38243 18955
rect 39221 18921 39255 18955
rect 40785 18921 40819 18955
rect 42809 18921 42843 18955
rect 46489 18921 46523 18955
rect 47501 18921 47535 18955
rect 51089 18921 51123 18955
rect 55505 18921 55539 18955
rect 26617 18853 26651 18887
rect 39129 18853 39163 18887
rect 30297 18785 30331 18819
rect 32781 18785 32815 18819
rect 32873 18785 32907 18819
rect 35817 18785 35851 18819
rect 40141 18785 40175 18819
rect 40509 18785 40543 18819
rect 41521 18785 41555 18819
rect 41797 18785 41831 18819
rect 43453 18785 43487 18819
rect 50537 18785 50571 18819
rect 52745 18785 52779 18819
rect 55781 18785 55815 18819
rect 21557 18717 21591 18751
rect 22017 18717 22051 18751
rect 22201 18717 22235 18751
rect 23121 18717 23155 18751
rect 23305 18717 23339 18751
rect 24041 18717 24075 18751
rect 25513 18717 25547 18751
rect 25605 18717 25639 18751
rect 29009 18717 29043 18751
rect 30389 18717 30423 18751
rect 31769 18717 31803 18751
rect 32045 18717 32079 18751
rect 32689 18717 32723 18751
rect 32965 18717 32999 18751
rect 35173 18717 35207 18751
rect 35357 18717 35391 18751
rect 36001 18717 36035 18751
rect 36185 18717 36219 18751
rect 36737 18717 36771 18751
rect 36921 18717 36955 18751
rect 38853 18717 38887 18751
rect 38991 18717 39025 18751
rect 39313 18717 39347 18751
rect 40601 18717 40635 18751
rect 41429 18717 41463 18751
rect 43177 18717 43211 18751
rect 46673 18717 46707 18751
rect 46949 18717 46983 18751
rect 47409 18717 47443 18751
rect 47593 18717 47627 18751
rect 50629 18717 50663 18751
rect 50721 18717 50755 18751
rect 52101 18717 52135 18751
rect 52377 18717 52411 18751
rect 53665 18717 53699 18751
rect 55689 18717 55723 18751
rect 58081 18717 58115 18751
rect 23213 18649 23247 18683
rect 26249 18649 26283 18683
rect 26433 18649 26467 18683
rect 31953 18649 31987 18683
rect 37841 18649 37875 18683
rect 38025 18649 38059 18683
rect 46857 18649 46891 18683
rect 54401 18649 54435 18683
rect 56609 18649 56643 18683
rect 24593 18581 24627 18615
rect 25789 18581 25823 18615
rect 36737 18581 36771 18615
rect 43269 18581 43303 18615
rect 44097 18581 44131 18615
rect 45293 18581 45327 18615
rect 45937 18581 45971 18615
rect 48053 18581 48087 18615
rect 48697 18581 48731 18615
rect 49249 18581 49283 18615
rect 49801 18581 49835 18615
rect 56149 18581 56183 18615
rect 57253 18581 57287 18615
rect 58265 18581 58299 18615
rect 24501 18377 24535 18411
rect 24685 18377 24719 18411
rect 25789 18377 25823 18411
rect 26617 18377 26651 18411
rect 28365 18377 28399 18411
rect 30021 18377 30055 18411
rect 35633 18377 35667 18411
rect 35817 18377 35851 18411
rect 38301 18377 38335 18411
rect 39773 18377 39807 18411
rect 41245 18377 41279 18411
rect 44097 18377 44131 18411
rect 53389 18377 53423 18411
rect 55137 18377 55171 18411
rect 24869 18309 24903 18343
rect 27261 18309 27295 18343
rect 37473 18309 37507 18343
rect 46397 18309 46431 18343
rect 53757 18309 53791 18343
rect 55689 18309 55723 18343
rect 1593 18241 1627 18275
rect 22017 18241 22051 18275
rect 24777 18241 24811 18275
rect 25053 18241 25087 18275
rect 25513 18241 25547 18275
rect 25605 18241 25639 18275
rect 26249 18241 26283 18275
rect 27169 18241 27203 18275
rect 27997 18241 28031 18275
rect 28181 18241 28215 18275
rect 29561 18241 29595 18275
rect 29837 18241 29871 18275
rect 30481 18241 30515 18275
rect 31125 18241 31159 18275
rect 32873 18241 32907 18275
rect 32965 18241 32999 18275
rect 33149 18241 33183 18275
rect 35758 18241 35792 18275
rect 36185 18241 36219 18275
rect 37749 18241 37783 18275
rect 38209 18241 38243 18275
rect 38393 18241 38427 18275
rect 39313 18241 39347 18275
rect 39589 18241 39623 18275
rect 41245 18241 41279 18275
rect 41429 18241 41463 18275
rect 42809 18241 42843 18275
rect 43361 18241 43395 18275
rect 43821 18241 43855 18275
rect 44741 18241 44775 18275
rect 45661 18241 45695 18275
rect 45845 18241 45879 18275
rect 45937 18241 45971 18275
rect 46213 18241 46247 18275
rect 48329 18241 48363 18275
rect 48513 18241 48547 18275
rect 48973 18241 49007 18275
rect 49157 18241 49191 18275
rect 50169 18241 50203 18275
rect 50353 18241 50387 18275
rect 53573 18241 53607 18275
rect 53665 18241 53699 18275
rect 53941 18241 53975 18275
rect 55045 18241 55079 18275
rect 55781 18241 55815 18275
rect 55965 18241 55999 18275
rect 57069 18241 57103 18275
rect 58081 18241 58115 18275
rect 22293 18173 22327 18207
rect 24041 18173 24075 18207
rect 25789 18173 25823 18207
rect 26341 18173 26375 18207
rect 27905 18173 27939 18207
rect 28089 18173 28123 18207
rect 30573 18173 30607 18207
rect 36277 18173 36311 18207
rect 37473 18173 37507 18207
rect 39405 18173 39439 18207
rect 44097 18173 44131 18207
rect 44649 18173 44683 18207
rect 46029 18173 46063 18207
rect 46857 18173 46891 18207
rect 49065 18173 49099 18207
rect 29653 18105 29687 18139
rect 29745 18105 29779 18139
rect 33149 18105 33183 18139
rect 45109 18105 45143 18139
rect 48329 18105 48363 18139
rect 50905 18105 50939 18139
rect 56517 18105 56551 18139
rect 1777 18037 1811 18071
rect 26249 18037 26283 18071
rect 36829 18037 36863 18071
rect 37657 18037 37691 18071
rect 39313 18037 39347 18071
rect 43913 18037 43947 18071
rect 48053 18037 48087 18071
rect 49985 18037 50019 18071
rect 51457 18037 51491 18071
rect 51917 18037 51951 18071
rect 54401 18037 54435 18071
rect 23305 17833 23339 17867
rect 24593 17833 24627 17867
rect 26341 17833 26375 17867
rect 28089 17833 28123 17867
rect 29009 17833 29043 17867
rect 33793 17833 33827 17867
rect 35265 17833 35299 17867
rect 36829 17833 36863 17867
rect 39037 17833 39071 17867
rect 39221 17833 39255 17867
rect 45201 17833 45235 17867
rect 48421 17833 48455 17867
rect 48605 17833 48639 17867
rect 50997 17833 51031 17867
rect 51825 17833 51859 17867
rect 53205 17833 53239 17867
rect 53849 17833 53883 17867
rect 54217 17833 54251 17867
rect 55505 17833 55539 17867
rect 57805 17833 57839 17867
rect 1593 17765 1627 17799
rect 23949 17765 23983 17799
rect 31309 17765 31343 17799
rect 43913 17765 43947 17799
rect 47593 17765 47627 17799
rect 49617 17765 49651 17799
rect 52101 17765 52135 17799
rect 53389 17765 53423 17799
rect 24041 17697 24075 17731
rect 24777 17697 24811 17731
rect 24869 17697 24903 17731
rect 27537 17697 27571 17731
rect 29101 17697 29135 17731
rect 31033 17697 31067 17731
rect 33885 17697 33919 17731
rect 34897 17697 34931 17731
rect 37105 17697 37139 17731
rect 43545 17697 43579 17731
rect 44465 17697 44499 17731
rect 49801 17697 49835 17731
rect 52193 17697 52227 17731
rect 52285 17697 52319 17731
rect 55965 17697 55999 17731
rect 56149 17697 56183 17731
rect 23765 17629 23799 17663
rect 23857 17629 23891 17663
rect 24961 17629 24995 17663
rect 25053 17629 25087 17663
rect 27261 17629 27295 17663
rect 27353 17629 27387 17663
rect 27997 17629 28031 17663
rect 28089 17629 28123 17663
rect 28365 17629 28399 17663
rect 29193 17629 29227 17663
rect 30941 17629 30975 17663
rect 32413 17629 32447 17663
rect 32597 17629 32631 17663
rect 32781 17629 32815 17663
rect 33057 17629 33091 17663
rect 33149 17629 33183 17663
rect 33609 17629 33643 17663
rect 33701 17629 33735 17663
rect 35081 17629 35115 17663
rect 37013 17629 37047 17663
rect 37197 17629 37231 17663
rect 37289 17629 37323 17663
rect 37473 17629 37507 17663
rect 37933 17629 37967 17663
rect 43269 17629 43303 17663
rect 43453 17629 43487 17663
rect 43637 17629 43671 17663
rect 43729 17629 43763 17663
rect 44557 17629 44591 17663
rect 45385 17629 45419 17663
rect 45477 17629 45511 17663
rect 45661 17629 45695 17663
rect 45753 17629 45787 17663
rect 46397 17629 46431 17663
rect 46489 17629 46523 17663
rect 46857 17629 46891 17663
rect 49525 17629 49559 17663
rect 50353 17629 50387 17663
rect 50537 17629 50571 17663
rect 50629 17629 50663 17663
rect 50721 17629 50755 17663
rect 52009 17629 52043 17663
rect 52469 17629 52503 17663
rect 53849 17629 53883 17663
rect 54033 17629 54067 17663
rect 55873 17629 55907 17663
rect 26157 17561 26191 17595
rect 26362 17561 26396 17595
rect 38025 17561 38059 17595
rect 38853 17561 38887 17595
rect 46673 17561 46707 17595
rect 46763 17561 46797 17595
rect 48237 17561 48271 17595
rect 53021 17561 53055 17595
rect 25605 17493 25639 17527
rect 26525 17493 26559 17527
rect 27537 17493 27571 17527
rect 28181 17493 28215 17527
rect 28825 17493 28859 17527
rect 39053 17493 39087 17527
rect 40601 17493 40635 17527
rect 42717 17493 42751 17527
rect 47041 17493 47075 17527
rect 48437 17493 48471 17527
rect 49801 17493 49835 17527
rect 53221 17493 53255 17527
rect 54677 17493 54711 17527
rect 56701 17493 56735 17527
rect 57345 17493 57379 17527
rect 22477 17289 22511 17323
rect 24961 17289 24995 17323
rect 25605 17289 25639 17323
rect 31217 17289 31251 17323
rect 32689 17289 32723 17323
rect 34069 17289 34103 17323
rect 35265 17289 35299 17323
rect 35725 17289 35759 17323
rect 37473 17289 37507 17323
rect 38853 17289 38887 17323
rect 40233 17289 40267 17323
rect 40877 17289 40911 17323
rect 42993 17289 43027 17323
rect 43821 17289 43855 17323
rect 46121 17289 46155 17323
rect 46765 17289 46799 17323
rect 50353 17289 50387 17323
rect 51549 17289 51583 17323
rect 53941 17289 53975 17323
rect 54493 17289 54527 17323
rect 56425 17289 56459 17323
rect 57437 17289 57471 17323
rect 27813 17221 27847 17255
rect 34805 17221 34839 17255
rect 36093 17221 36127 17255
rect 40693 17221 40727 17255
rect 47777 17221 47811 17255
rect 54677 17221 54711 17255
rect 22569 17153 22603 17187
rect 24593 17153 24627 17187
rect 25421 17153 25455 17187
rect 26341 17153 26375 17187
rect 26525 17153 26559 17187
rect 27997 17153 28031 17187
rect 29193 17153 29227 17187
rect 29285 17153 29319 17187
rect 29469 17153 29503 17187
rect 29929 17153 29963 17187
rect 30573 17153 30607 17187
rect 30757 17153 30791 17187
rect 30849 17153 30883 17187
rect 30941 17153 30975 17187
rect 32505 17153 32539 17187
rect 33701 17153 33735 17187
rect 33885 17153 33919 17187
rect 34897 17153 34931 17187
rect 36185 17153 36219 17187
rect 37749 17153 37783 17187
rect 38761 17153 38795 17187
rect 39037 17153 39071 17187
rect 39957 17153 39991 17187
rect 40141 17153 40175 17187
rect 40233 17153 40267 17187
rect 42717 17153 42751 17187
rect 43453 17153 43487 17187
rect 43637 17153 43671 17187
rect 44649 17153 44683 17187
rect 44833 17153 44867 17187
rect 45937 17153 45971 17187
rect 46121 17153 46155 17187
rect 46949 17153 46983 17187
rect 47133 17153 47167 17187
rect 48973 17153 49007 17187
rect 49525 17153 49559 17187
rect 50445 17153 50479 17187
rect 50997 17153 51031 17187
rect 51181 17153 51215 17187
rect 51273 17153 51307 17187
rect 51365 17153 51399 17187
rect 52009 17153 52043 17187
rect 53297 17153 53331 17187
rect 53849 17153 53883 17187
rect 54033 17153 54067 17187
rect 54861 17153 54895 17187
rect 55873 17153 55907 17187
rect 56149 17153 56183 17187
rect 56241 17153 56275 17187
rect 24685 17085 24719 17119
rect 32321 17085 32355 17119
rect 34621 17085 34655 17119
rect 36277 17085 36311 17119
rect 37473 17085 37507 17119
rect 42993 17085 43027 17119
rect 47225 17085 47259 17119
rect 49249 17085 49283 17119
rect 49709 17085 49743 17119
rect 52101 17085 52135 17119
rect 52285 17085 52319 17119
rect 56885 17085 56919 17119
rect 58081 17085 58115 17119
rect 39037 17017 39071 17051
rect 42073 17017 42107 17051
rect 44741 17017 44775 17051
rect 52193 17017 52227 17051
rect 55413 17017 55447 17051
rect 23857 16949 23891 16983
rect 24777 16949 24811 16983
rect 26525 16949 26559 16983
rect 27629 16949 27663 16983
rect 28641 16949 28675 16983
rect 29469 16949 29503 16983
rect 37657 16949 37691 16983
rect 40877 16949 40911 16983
rect 41061 16949 41095 16983
rect 42809 16949 42843 16983
rect 43453 16949 43487 16983
rect 45293 16949 45327 16983
rect 53021 16949 53055 16983
rect 55965 16949 55999 16983
rect 24041 16745 24075 16779
rect 29009 16745 29043 16779
rect 31217 16745 31251 16779
rect 40509 16745 40543 16779
rect 44097 16745 44131 16779
rect 52469 16745 52503 16779
rect 52837 16745 52871 16779
rect 53757 16745 53791 16779
rect 54493 16745 54527 16779
rect 56057 16745 56091 16779
rect 56609 16745 56643 16779
rect 26525 16677 26559 16711
rect 27905 16677 27939 16711
rect 29193 16677 29227 16711
rect 36737 16677 36771 16711
rect 37105 16677 37139 16711
rect 48973 16677 49007 16711
rect 22293 16609 22327 16643
rect 22569 16609 22603 16643
rect 26249 16609 26283 16643
rect 27629 16609 27663 16643
rect 29929 16609 29963 16643
rect 33333 16609 33367 16643
rect 37013 16609 37047 16643
rect 38393 16609 38427 16643
rect 39313 16609 39347 16643
rect 48145 16609 48179 16643
rect 52377 16609 52411 16643
rect 56517 16609 56551 16643
rect 56701 16609 56735 16643
rect 26157 16541 26191 16575
rect 27537 16541 27571 16575
rect 30021 16541 30055 16575
rect 30297 16541 30331 16575
rect 31125 16541 31159 16575
rect 31309 16541 31343 16575
rect 31953 16541 31987 16575
rect 33977 16541 34011 16575
rect 34161 16541 34195 16575
rect 36921 16541 36955 16575
rect 37197 16541 37231 16575
rect 37381 16541 37415 16575
rect 38301 16541 38335 16575
rect 39129 16541 39163 16575
rect 39497 16541 39531 16575
rect 40049 16541 40083 16575
rect 40141 16541 40175 16575
rect 40325 16541 40359 16575
rect 41521 16541 41555 16575
rect 41981 16541 42015 16575
rect 45845 16541 45879 16575
rect 46121 16541 46155 16575
rect 46213 16541 46247 16575
rect 46489 16541 46523 16575
rect 46673 16541 46707 16575
rect 47777 16541 47811 16575
rect 47961 16541 47995 16575
rect 48237 16541 48271 16575
rect 48513 16541 48547 16575
rect 49157 16541 49191 16575
rect 50537 16541 50571 16575
rect 50721 16541 50755 16575
rect 51365 16541 51399 16575
rect 51457 16541 51491 16575
rect 51733 16541 51767 16575
rect 52653 16541 52687 16575
rect 53297 16541 53331 16575
rect 53573 16541 53607 16575
rect 54677 16541 54711 16575
rect 54769 16541 54803 16575
rect 55505 16541 55539 16575
rect 55597 16541 55631 16575
rect 55781 16541 55815 16575
rect 55873 16541 55907 16575
rect 56793 16541 56827 16575
rect 29055 16507 29089 16541
rect 24685 16473 24719 16507
rect 28825 16473 28859 16507
rect 33241 16473 33275 16507
rect 39221 16473 39255 16507
rect 43821 16473 43855 16507
rect 45385 16473 45419 16507
rect 49341 16473 49375 16507
rect 50629 16473 50663 16507
rect 51549 16473 51583 16507
rect 54493 16473 54527 16507
rect 30297 16405 30331 16439
rect 31861 16405 31895 16439
rect 32781 16405 32815 16439
rect 33149 16405 33183 16439
rect 34161 16405 34195 16439
rect 37841 16405 37875 16439
rect 38209 16405 38243 16439
rect 39405 16405 39439 16439
rect 51181 16405 51215 16439
rect 53389 16405 53423 16439
rect 57253 16405 57287 16439
rect 57897 16405 57931 16439
rect 23765 16201 23799 16235
rect 25513 16201 25547 16235
rect 26617 16201 26651 16235
rect 29193 16201 29227 16235
rect 30113 16201 30147 16235
rect 31585 16201 31619 16235
rect 33241 16201 33275 16235
rect 34345 16201 34379 16235
rect 34713 16201 34747 16235
rect 36829 16201 36863 16235
rect 38117 16201 38151 16235
rect 40325 16201 40359 16235
rect 40693 16201 40727 16235
rect 41153 16201 41187 16235
rect 41797 16201 41831 16235
rect 42809 16201 42843 16235
rect 44741 16201 44775 16235
rect 46213 16201 46247 16235
rect 46765 16201 46799 16235
rect 48513 16201 48547 16235
rect 49525 16201 49559 16235
rect 50169 16201 50203 16235
rect 51733 16201 51767 16235
rect 53665 16201 53699 16235
rect 55137 16201 55171 16235
rect 56057 16201 56091 16235
rect 22293 16133 22327 16167
rect 27629 16133 27663 16167
rect 34805 16133 34839 16167
rect 42993 16133 43027 16167
rect 44373 16133 44407 16167
rect 51273 16133 51307 16167
rect 22017 16065 22051 16099
rect 24593 16065 24627 16099
rect 26433 16065 26467 16099
rect 27445 16065 27479 16099
rect 29745 16065 29779 16099
rect 29929 16065 29963 16099
rect 31033 16065 31067 16099
rect 31125 16065 31159 16099
rect 31309 16065 31343 16099
rect 31401 16065 31435 16099
rect 32873 16065 32907 16099
rect 32965 16065 32999 16099
rect 35725 16065 35759 16099
rect 36737 16065 36771 16099
rect 36921 16065 36955 16099
rect 38025 16065 38059 16099
rect 38209 16065 38243 16099
rect 40233 16065 40267 16099
rect 40509 16065 40543 16099
rect 41521 16065 41555 16099
rect 41613 16065 41647 16099
rect 42717 16065 42751 16099
rect 43545 16065 43579 16099
rect 43729 16065 43763 16099
rect 44557 16065 44591 16099
rect 45569 16065 45603 16099
rect 45752 16065 45786 16099
rect 45937 16065 45971 16099
rect 46121 16065 46155 16099
rect 46765 16065 46799 16099
rect 46949 16065 46983 16099
rect 47777 16065 47811 16099
rect 47961 16065 47995 16099
rect 48697 16065 48731 16099
rect 48881 16065 48915 16099
rect 50353 16065 50387 16099
rect 50629 16065 50663 16099
rect 50813 16065 50847 16099
rect 51549 16065 51583 16099
rect 52193 16065 52227 16099
rect 53849 16065 53883 16099
rect 54033 16065 54067 16099
rect 54861 16065 54895 16099
rect 55965 16065 55999 16099
rect 56149 16065 56183 16099
rect 24685 15997 24719 16031
rect 24961 15997 24995 16031
rect 26157 15997 26191 16031
rect 26249 15997 26283 16031
rect 26341 15997 26375 16031
rect 27169 15997 27203 16031
rect 32781 15997 32815 16031
rect 33057 15997 33091 16031
rect 34989 15997 35023 16031
rect 35633 15997 35667 16031
rect 45845 15997 45879 16031
rect 48789 15997 48823 16031
rect 48973 15997 49007 16031
rect 51365 15997 51399 16031
rect 53941 15997 53975 16031
rect 54125 15997 54159 16031
rect 28181 15929 28215 15963
rect 36093 15929 36127 15963
rect 43637 15929 43671 15963
rect 47961 15929 47995 15963
rect 50445 15929 50479 15963
rect 50537 15929 50571 15963
rect 58081 15929 58115 15963
rect 27261 15861 27295 15895
rect 28641 15861 28675 15895
rect 29745 15861 29779 15895
rect 38761 15861 38795 15895
rect 42993 15861 43027 15895
rect 51273 15861 51307 15895
rect 53021 15861 53055 15895
rect 56609 15861 56643 15895
rect 57161 15861 57195 15895
rect 25421 15657 25455 15691
rect 26617 15657 26651 15691
rect 31033 15657 31067 15691
rect 32965 15657 32999 15691
rect 35633 15657 35667 15691
rect 36093 15657 36127 15691
rect 37657 15657 37691 15691
rect 38485 15657 38519 15691
rect 41981 15657 42015 15691
rect 46121 15657 46155 15691
rect 50813 15657 50847 15691
rect 51917 15657 51951 15691
rect 54953 15657 54987 15691
rect 57529 15657 57563 15691
rect 24777 15589 24811 15623
rect 27905 15589 27939 15623
rect 27997 15589 28031 15623
rect 32505 15589 32539 15623
rect 42533 15589 42567 15623
rect 43361 15589 43395 15623
rect 44281 15589 44315 15623
rect 46489 15589 46523 15623
rect 21833 15521 21867 15555
rect 29837 15521 29871 15555
rect 30297 15521 30331 15555
rect 35173 15521 35207 15555
rect 39037 15521 39071 15555
rect 42993 15521 43027 15555
rect 45385 15521 45419 15555
rect 46397 15521 46431 15555
rect 47409 15521 47443 15555
rect 47501 15521 47535 15555
rect 47685 15521 47719 15555
rect 51273 15521 51307 15555
rect 52377 15521 52411 15555
rect 58081 15521 58115 15555
rect 22477 15453 22511 15487
rect 22661 15453 22695 15487
rect 23581 15453 23615 15487
rect 24593 15453 24627 15487
rect 26065 15453 26099 15487
rect 26157 15453 26191 15487
rect 26341 15453 26375 15487
rect 26433 15453 26467 15487
rect 28733 15453 28767 15487
rect 28825 15453 28859 15487
rect 29009 15453 29043 15487
rect 29101 15453 29135 15487
rect 29929 15453 29963 15487
rect 31309 15453 31343 15487
rect 32137 15453 32171 15487
rect 32965 15453 32999 15487
rect 33241 15453 33275 15487
rect 34897 15453 34931 15487
rect 35081 15453 35115 15487
rect 35265 15453 35299 15487
rect 35449 15453 35483 15487
rect 36277 15453 36311 15487
rect 36645 15453 36679 15487
rect 37197 15453 37231 15487
rect 37657 15453 37691 15487
rect 37933 15453 37967 15487
rect 43177 15453 43211 15487
rect 45201 15453 45235 15487
rect 45569 15453 45603 15487
rect 46305 15453 46339 15487
rect 46581 15453 46615 15487
rect 47593 15453 47627 15487
rect 50353 15453 50387 15487
rect 50629 15453 50663 15487
rect 52101 15453 52135 15487
rect 52285 15453 52319 15487
rect 53021 15453 53055 15487
rect 53205 15453 53239 15487
rect 53297 15453 53331 15487
rect 55965 15453 55999 15487
rect 56977 15453 57011 15487
rect 27537 15385 27571 15419
rect 31033 15385 31067 15419
rect 32321 15385 32355 15419
rect 36369 15385 36403 15419
rect 36461 15385 36495 15419
rect 38945 15385 38979 15419
rect 44005 15385 44039 15419
rect 48329 15385 48363 15419
rect 48881 15385 48915 15419
rect 49433 15385 49467 15419
rect 49617 15385 49651 15419
rect 55597 15385 55631 15419
rect 22293 15317 22327 15351
rect 23397 15317 23431 15351
rect 28549 15317 28583 15351
rect 31217 15317 31251 15351
rect 33149 15317 33183 15351
rect 34345 15317 34379 15351
rect 37841 15317 37875 15351
rect 38853 15317 38887 15351
rect 40049 15317 40083 15351
rect 45293 15317 45327 15351
rect 45477 15317 45511 15351
rect 47869 15317 47903 15351
rect 49801 15317 49835 15351
rect 50445 15317 50479 15351
rect 52837 15317 52871 15351
rect 53757 15317 53791 15351
rect 54309 15317 54343 15351
rect 56425 15317 56459 15351
rect 23673 15113 23707 15147
rect 24041 15113 24075 15147
rect 24869 15113 24903 15147
rect 25789 15113 25823 15147
rect 28733 15113 28767 15147
rect 30389 15113 30423 15147
rect 36461 15113 36495 15147
rect 37841 15113 37875 15147
rect 38945 15113 38979 15147
rect 41705 15113 41739 15147
rect 43361 15113 43395 15147
rect 44649 15113 44683 15147
rect 47977 15113 48011 15147
rect 48145 15113 48179 15147
rect 53129 15113 53163 15147
rect 53297 15113 53331 15147
rect 53849 15113 53883 15147
rect 22845 15045 22879 15079
rect 26525 15045 26559 15079
rect 27261 15045 27295 15079
rect 31033 15045 31067 15079
rect 32873 15045 32907 15079
rect 34069 15045 34103 15079
rect 34713 15045 34747 15079
rect 46949 15045 46983 15079
rect 47777 15045 47811 15079
rect 51181 15045 51215 15079
rect 52377 15045 52411 15079
rect 52929 15045 52963 15079
rect 22477 14977 22511 15011
rect 25605 14977 25639 15011
rect 26249 14977 26283 15011
rect 26341 14977 26375 15011
rect 27445 14977 27479 15011
rect 27629 14977 27663 15011
rect 27721 14977 27755 15011
rect 28917 14977 28951 15011
rect 30021 14977 30055 15011
rect 30205 14977 30239 15011
rect 31622 14977 31656 15011
rect 31769 14977 31803 15011
rect 34529 14977 34563 15011
rect 34897 14977 34931 15011
rect 35357 14977 35391 15011
rect 35541 14977 35575 15011
rect 36369 14977 36403 15011
rect 36553 14977 36587 15011
rect 37473 14977 37507 15011
rect 39313 14977 39347 15011
rect 40693 14977 40727 15011
rect 40877 14977 40911 15011
rect 43545 14977 43579 15011
rect 43637 14977 43671 15011
rect 43729 14977 43763 15011
rect 44833 14977 44867 15011
rect 44925 14977 44959 15011
rect 45109 14977 45143 15011
rect 45661 14977 45695 15011
rect 45753 14977 45787 15011
rect 45937 14977 45971 15011
rect 46029 14977 46063 15011
rect 46765 14977 46799 15011
rect 48605 14977 48639 15011
rect 48789 14977 48823 15011
rect 48973 14977 49007 15011
rect 49065 14977 49099 15011
rect 49893 14977 49927 15011
rect 50214 14977 50248 15011
rect 50353 14977 50387 15011
rect 50905 14977 50939 15011
rect 51089 14977 51123 15011
rect 52101 14977 52135 15011
rect 52193 14977 52227 15011
rect 54033 14977 54067 15011
rect 54125 14977 54159 15011
rect 54309 14977 54343 15011
rect 54401 14977 54435 15011
rect 55229 14977 55263 15011
rect 55505 14977 55539 15011
rect 55689 14977 55723 15011
rect 56057 14977 56091 15011
rect 56609 14977 56643 15011
rect 56977 14977 57011 15011
rect 24133 14909 24167 14943
rect 24317 14909 24351 14943
rect 25421 14909 25455 14943
rect 29193 14909 29227 14943
rect 31401 14909 31435 14943
rect 32413 14909 32447 14943
rect 37565 14909 37599 14943
rect 39129 14909 39163 14943
rect 39221 14909 39255 14943
rect 39405 14909 39439 14943
rect 46213 14909 46247 14943
rect 48881 14909 48915 14943
rect 49709 14909 49743 14943
rect 49985 14909 50019 14943
rect 50077 14909 50111 14943
rect 26525 14841 26559 14875
rect 31493 14841 31527 14875
rect 35449 14841 35483 14875
rect 43913 14841 43947 14875
rect 45017 14841 45051 14875
rect 49249 14841 49283 14875
rect 52377 14841 52411 14875
rect 21373 14773 21407 14807
rect 28273 14773 28307 14807
rect 29101 14773 29135 14807
rect 33425 14773 33459 14807
rect 37473 14773 37507 14807
rect 38301 14773 38335 14807
rect 39957 14773 39991 14807
rect 42901 14773 42935 14807
rect 47133 14773 47167 14807
rect 47961 14773 47995 14807
rect 53113 14773 53147 14807
rect 58081 14773 58115 14807
rect 24593 14569 24627 14603
rect 26801 14569 26835 14603
rect 31861 14569 31895 14603
rect 32965 14569 32999 14603
rect 33425 14569 33459 14603
rect 35541 14569 35575 14603
rect 36553 14569 36587 14603
rect 36737 14569 36771 14603
rect 37933 14569 37967 14603
rect 38393 14569 38427 14603
rect 40601 14569 40635 14603
rect 41429 14569 41463 14603
rect 43729 14569 43763 14603
rect 44465 14569 44499 14603
rect 45661 14569 45695 14603
rect 46857 14569 46891 14603
rect 48053 14569 48087 14603
rect 48973 14569 49007 14603
rect 51181 14569 51215 14603
rect 52561 14569 52595 14603
rect 53021 14569 53055 14603
rect 54401 14569 54435 14603
rect 56241 14569 56275 14603
rect 57345 14569 57379 14603
rect 22569 14501 22603 14535
rect 42625 14501 42659 14535
rect 49801 14501 49835 14535
rect 50997 14501 51031 14535
rect 51089 14501 51123 14535
rect 23029 14433 23063 14467
rect 25145 14433 25179 14467
rect 27353 14433 27387 14467
rect 28365 14433 28399 14467
rect 37473 14433 37507 14467
rect 40417 14433 40451 14467
rect 42717 14433 42751 14467
rect 50813 14433 50847 14467
rect 52193 14433 52227 14467
rect 55597 14433 55631 14467
rect 22385 14365 22419 14399
rect 23305 14365 23339 14399
rect 27537 14365 27571 14399
rect 27813 14365 27847 14399
rect 31217 14365 31251 14399
rect 31401 14365 31435 14399
rect 31493 14365 31527 14399
rect 31585 14365 31619 14399
rect 32321 14365 32355 14399
rect 32505 14365 32539 14399
rect 32597 14365 32631 14399
rect 32735 14365 32769 14399
rect 33612 14343 33646 14377
rect 33701 14365 33735 14399
rect 33897 14365 33931 14399
rect 33987 14365 34021 14399
rect 34897 14365 34931 14399
rect 35081 14365 35115 14399
rect 35173 14365 35207 14399
rect 35265 14365 35299 14399
rect 37565 14365 37599 14399
rect 37749 14365 37783 14399
rect 38577 14365 38611 14399
rect 38853 14365 38887 14399
rect 39037 14365 39071 14399
rect 40325 14365 40359 14399
rect 41613 14365 41647 14399
rect 41889 14365 41923 14399
rect 42441 14365 42475 14399
rect 42533 14365 42567 14399
rect 42809 14365 42843 14399
rect 45891 14365 45925 14399
rect 46042 14365 46076 14399
rect 46142 14359 46176 14393
rect 46305 14365 46339 14399
rect 47041 14365 47075 14399
rect 47133 14365 47167 14399
rect 47409 14365 47443 14399
rect 47501 14365 47535 14399
rect 48237 14365 48271 14399
rect 48513 14365 48547 14399
rect 49157 14365 49191 14399
rect 49249 14365 49283 14399
rect 51273 14365 51307 14399
rect 51917 14365 51951 14399
rect 52101 14365 52135 14399
rect 52285 14365 52319 14399
rect 52377 14365 52411 14399
rect 53205 14365 53239 14399
rect 53297 14365 53331 14399
rect 53481 14365 53515 14399
rect 53573 14365 53607 14399
rect 54033 14365 54067 14399
rect 54217 14365 54251 14399
rect 55505 14365 55539 14399
rect 55689 14365 55723 14399
rect 24961 14297 24995 14331
rect 26525 14297 26559 14331
rect 27721 14297 27755 14331
rect 36093 14297 36127 14331
rect 36921 14297 36955 14331
rect 43545 14297 43579 14331
rect 47225 14297 47259 14331
rect 48973 14297 49007 14331
rect 24041 14229 24075 14263
rect 25053 14229 25087 14263
rect 25973 14229 26007 14263
rect 28917 14229 28951 14263
rect 36721 14229 36755 14263
rect 41797 14229 41831 14263
rect 43745 14229 43779 14263
rect 43913 14229 43947 14263
rect 48421 14229 48455 14263
rect 51365 14229 51399 14263
rect 54861 14229 54895 14263
rect 56701 14229 56735 14263
rect 57805 14229 57839 14263
rect 28733 14025 28767 14059
rect 29377 14025 29411 14059
rect 30855 14025 30889 14059
rect 32321 14025 32355 14059
rect 34529 14025 34563 14059
rect 35633 14025 35667 14059
rect 37473 14025 37507 14059
rect 38577 14025 38611 14059
rect 38761 14025 38795 14059
rect 41613 14025 41647 14059
rect 43637 14025 43671 14059
rect 45477 14025 45511 14059
rect 47225 14025 47259 14059
rect 50629 14025 50663 14059
rect 51181 14025 51215 14059
rect 52285 14025 52319 14059
rect 53573 14025 53607 14059
rect 54493 14025 54527 14059
rect 55137 14025 55171 14059
rect 58081 14025 58115 14059
rect 26249 13957 26283 13991
rect 30757 13957 30791 13991
rect 34897 13957 34931 13991
rect 36001 13957 36035 13991
rect 43453 13957 43487 13991
rect 53205 13957 53239 13991
rect 55689 13957 55723 13991
rect 24961 13889 24995 13923
rect 25421 13889 25455 13923
rect 25605 13889 25639 13923
rect 26341 13889 26375 13923
rect 26617 13889 26651 13923
rect 27813 13889 27847 13923
rect 27997 13889 28031 13923
rect 28089 13889 28123 13923
rect 28641 13889 28675 13923
rect 28825 13889 28859 13923
rect 29377 13889 29411 13923
rect 29561 13889 29595 13923
rect 29653 13889 29687 13923
rect 29929 13889 29963 13923
rect 30941 13889 30975 13923
rect 31033 13889 31067 13923
rect 32505 13889 32539 13923
rect 32689 13889 32723 13923
rect 32781 13889 32815 13923
rect 33241 13889 33275 13923
rect 33425 13889 33459 13923
rect 33517 13889 33551 13923
rect 33645 13889 33679 13923
rect 34437 13889 34471 13923
rect 34713 13889 34747 13923
rect 35817 13889 35851 13923
rect 35909 13889 35943 13923
rect 36185 13889 36219 13923
rect 36737 13889 36771 13923
rect 36921 13889 36955 13923
rect 37657 13889 37691 13923
rect 38758 13889 38792 13923
rect 39221 13889 39255 13923
rect 39865 13889 39899 13923
rect 40049 13889 40083 13923
rect 40509 13889 40543 13923
rect 41429 13889 41463 13923
rect 42717 13889 42751 13923
rect 43269 13889 43303 13923
rect 44741 13889 44775 13923
rect 45385 13889 45419 13923
rect 45569 13889 45603 13923
rect 46489 13889 46523 13923
rect 46673 13889 46707 13923
rect 46857 13889 46891 13923
rect 47041 13889 47075 13923
rect 48789 13889 48823 13923
rect 48973 13889 49007 13923
rect 51089 13889 51123 13923
rect 51273 13889 51307 13923
rect 52193 13889 52227 13923
rect 52377 13889 52411 13923
rect 53113 13889 53147 13923
rect 53389 13889 53423 13923
rect 54217 13889 54251 13923
rect 54585 13889 54619 13923
rect 55781 13889 55815 13923
rect 56057 13889 56091 13923
rect 56701 13889 56735 13923
rect 56793 13889 56827 13923
rect 24225 13821 24259 13855
rect 27629 13821 27663 13855
rect 27905 13821 27939 13855
rect 29837 13821 29871 13855
rect 33333 13821 33367 13855
rect 36829 13821 36863 13855
rect 37841 13821 37875 13855
rect 39957 13821 39991 13855
rect 40969 13821 41003 13855
rect 46765 13821 46799 13855
rect 47777 13821 47811 13855
rect 49157 13821 49191 13855
rect 50169 13821 50203 13855
rect 50261 13821 50295 13855
rect 50353 13821 50387 13855
rect 50445 13821 50479 13855
rect 54033 13821 54067 13855
rect 24777 13753 24811 13787
rect 25697 13685 25731 13719
rect 39129 13685 39163 13719
rect 40601 13685 40635 13719
rect 44649 13685 44683 13719
rect 24961 13481 24995 13515
rect 25697 13481 25731 13515
rect 26065 13481 26099 13515
rect 31309 13481 31343 13515
rect 32321 13481 32355 13515
rect 33701 13481 33735 13515
rect 36093 13481 36127 13515
rect 37473 13481 37507 13515
rect 39221 13481 39255 13515
rect 40049 13481 40083 13515
rect 43085 13481 43119 13515
rect 44281 13481 44315 13515
rect 46397 13481 46431 13515
rect 47317 13481 47351 13515
rect 48697 13481 48731 13515
rect 52193 13481 52227 13515
rect 54677 13481 54711 13515
rect 56609 13481 56643 13515
rect 53665 13413 53699 13447
rect 54493 13413 54527 13447
rect 55505 13413 55539 13447
rect 30113 13345 30147 13379
rect 34345 13345 34379 13379
rect 37381 13345 37415 13379
rect 37565 13345 37599 13379
rect 40509 13345 40543 13379
rect 40693 13345 40727 13379
rect 42533 13345 42567 13379
rect 25881 13277 25915 13311
rect 26157 13277 26191 13311
rect 26893 13277 26927 13311
rect 27813 13277 27847 13311
rect 27997 13277 28031 13311
rect 28641 13277 28675 13311
rect 28733 13277 28767 13311
rect 28917 13277 28951 13311
rect 29009 13277 29043 13311
rect 29193 13277 29227 13311
rect 29929 13277 29963 13311
rect 30665 13277 30699 13311
rect 30849 13277 30883 13311
rect 30941 13277 30975 13311
rect 31033 13277 31067 13311
rect 31861 13277 31895 13311
rect 33241 13277 33275 13311
rect 33882 13277 33916 13311
rect 34253 13277 34287 13311
rect 35449 13277 35483 13311
rect 37289 13277 37323 13311
rect 38025 13277 38059 13311
rect 38209 13277 38243 13311
rect 41981 13277 42015 13311
rect 42349 13277 42383 13311
rect 42993 13277 43027 13311
rect 43177 13277 43211 13311
rect 43637 13277 43671 13311
rect 43785 13277 43819 13311
rect 44005 13277 44039 13311
rect 44143 13277 44177 13311
rect 45753 13277 45787 13311
rect 45916 13277 45950 13311
rect 46016 13277 46050 13311
rect 46121 13277 46155 13311
rect 47501 13277 47535 13311
rect 47593 13277 47627 13311
rect 47777 13277 47811 13311
rect 47869 13277 47903 13311
rect 49617 13277 49651 13311
rect 50353 13277 50387 13311
rect 50445 13277 50479 13311
rect 50629 13277 50663 13311
rect 51273 13277 51307 13311
rect 51457 13277 51491 13311
rect 51733 13277 51767 13311
rect 53573 13277 53607 13311
rect 55780 13255 55814 13289
rect 55873 13277 55907 13311
rect 55965 13277 55999 13311
rect 56149 13277 56183 13311
rect 58081 13277 58115 13311
rect 24869 13209 24903 13243
rect 26985 13209 27019 13243
rect 29745 13209 29779 13243
rect 36645 13209 36679 13243
rect 41245 13209 41279 13243
rect 43913 13209 43947 13243
rect 48329 13209 48363 13243
rect 48513 13209 48547 13243
rect 50813 13209 50847 13243
rect 54217 13209 54251 13243
rect 24041 13141 24075 13175
rect 27905 13141 27939 13175
rect 33885 13141 33919 13175
rect 34989 13141 35023 13175
rect 38117 13141 38151 13175
rect 38669 13141 38703 13175
rect 40417 13141 40451 13175
rect 42349 13141 42383 13175
rect 45201 13141 45235 13175
rect 49433 13141 49467 13175
rect 51641 13141 51675 13175
rect 52745 13141 52779 13175
rect 57161 13141 57195 13175
rect 58265 13141 58299 13175
rect 25881 12937 25915 12971
rect 28457 12937 28491 12971
rect 29101 12937 29135 12971
rect 31309 12937 31343 12971
rect 33333 12937 33367 12971
rect 34253 12937 34287 12971
rect 35725 12937 35759 12971
rect 36185 12937 36219 12971
rect 40969 12937 41003 12971
rect 42717 12937 42751 12971
rect 43085 12937 43119 12971
rect 45201 12937 45235 12971
rect 46305 12937 46339 12971
rect 47869 12937 47903 12971
rect 50537 12937 50571 12971
rect 24961 12869 24995 12903
rect 43729 12869 43763 12903
rect 44373 12869 44407 12903
rect 49341 12869 49375 12903
rect 51365 12869 51399 12903
rect 58081 12869 58115 12903
rect 23765 12801 23799 12835
rect 24317 12801 24351 12835
rect 24409 12801 24443 12835
rect 25145 12801 25179 12835
rect 25329 12801 25363 12835
rect 26065 12801 26099 12835
rect 26249 12801 26283 12835
rect 26525 12801 26559 12835
rect 27169 12801 27203 12835
rect 27445 12801 27479 12835
rect 27721 12801 27755 12835
rect 27905 12801 27939 12835
rect 29009 12801 29043 12835
rect 29193 12801 29227 12835
rect 29653 12801 29687 12835
rect 29837 12801 29871 12835
rect 31125 12801 31159 12835
rect 32689 12801 32723 12835
rect 33517 12801 33551 12835
rect 33609 12801 33643 12835
rect 33793 12801 33827 12835
rect 34989 12801 35023 12835
rect 35173 12801 35207 12835
rect 35541 12801 35575 12835
rect 36369 12801 36403 12835
rect 36553 12801 36587 12835
rect 36645 12801 36679 12835
rect 37565 12801 37599 12835
rect 38025 12801 38059 12835
rect 38209 12801 38243 12835
rect 38761 12801 38795 12835
rect 39037 12801 39071 12835
rect 41797 12801 41831 12835
rect 42901 12801 42935 12835
rect 43177 12801 43211 12835
rect 43821 12801 43855 12835
rect 45753 12801 45787 12835
rect 46949 12801 46983 12835
rect 47041 12801 47075 12835
rect 48053 12801 48087 12835
rect 48973 12801 49007 12835
rect 49121 12801 49155 12835
rect 49249 12801 49283 12835
rect 49438 12801 49472 12835
rect 50629 12801 50663 12835
rect 50813 12801 50847 12835
rect 52193 12801 52227 12835
rect 52377 12801 52411 12835
rect 52929 12801 52963 12835
rect 53205 12801 53239 12835
rect 54677 12801 54711 12835
rect 54861 12801 54895 12835
rect 55045 12801 55079 12835
rect 55505 12801 55539 12835
rect 25421 12733 25455 12767
rect 26341 12733 26375 12767
rect 27629 12733 27663 12767
rect 30849 12733 30883 12767
rect 32505 12733 32539 12767
rect 32597 12733 32631 12767
rect 32781 12733 32815 12767
rect 35265 12733 35299 12767
rect 35357 12733 35391 12767
rect 38945 12733 38979 12767
rect 40509 12733 40543 12767
rect 46029 12733 46063 12767
rect 46765 12733 46799 12767
rect 55781 12733 55815 12767
rect 26157 12665 26191 12699
rect 32321 12665 32355 12699
rect 38209 12665 38243 12699
rect 39221 12665 39255 12699
rect 40233 12665 40267 12699
rect 44557 12665 44591 12699
rect 53849 12665 53883 12699
rect 56885 12665 56919 12699
rect 29745 12597 29779 12631
rect 30941 12597 30975 12631
rect 33793 12597 33827 12631
rect 39037 12597 39071 12631
rect 40049 12597 40083 12631
rect 41981 12597 42015 12631
rect 46121 12597 46155 12631
rect 46857 12597 46891 12631
rect 49617 12597 49651 12631
rect 52377 12597 52411 12631
rect 53021 12597 53055 12631
rect 53389 12597 53423 12631
rect 55597 12597 55631 12631
rect 55689 12597 55723 12631
rect 56333 12597 56367 12631
rect 57437 12597 57471 12631
rect 24593 12393 24627 12427
rect 26065 12393 26099 12427
rect 27169 12393 27203 12427
rect 32321 12393 32355 12427
rect 33149 12393 33183 12427
rect 36737 12393 36771 12427
rect 37473 12393 37507 12427
rect 39313 12393 39347 12427
rect 40601 12393 40635 12427
rect 42165 12393 42199 12427
rect 43637 12393 43671 12427
rect 46397 12393 46431 12427
rect 49525 12393 49559 12427
rect 52929 12393 52963 12427
rect 53573 12393 53607 12427
rect 54401 12393 54435 12427
rect 56701 12393 56735 12427
rect 25513 12325 25547 12359
rect 40233 12325 40267 12359
rect 45201 12325 45235 12359
rect 47501 12325 47535 12359
rect 52653 12325 52687 12359
rect 53389 12325 53423 12359
rect 55505 12325 55539 12359
rect 27353 12257 27387 12291
rect 27445 12257 27479 12291
rect 27629 12257 27663 12291
rect 30573 12257 30607 12291
rect 33333 12257 33367 12291
rect 37841 12257 37875 12291
rect 50721 12257 50755 12291
rect 50813 12257 50847 12291
rect 51549 12257 51583 12291
rect 56057 12257 56091 12291
rect 27537 12189 27571 12223
rect 28549 12189 28583 12223
rect 28733 12189 28767 12223
rect 28825 12189 28859 12223
rect 28917 12189 28951 12223
rect 29009 12189 29043 12223
rect 30297 12189 30331 12223
rect 30481 12189 30515 12223
rect 30665 12189 30699 12223
rect 30849 12189 30883 12223
rect 31953 12189 31987 12223
rect 33425 12189 33459 12223
rect 33701 12189 33735 12223
rect 34897 12189 34931 12223
rect 35633 12189 35667 12223
rect 35817 12189 35851 12223
rect 36277 12189 36311 12223
rect 36553 12189 36587 12223
rect 37657 12189 37691 12223
rect 37933 12189 37967 12223
rect 38025 12189 38059 12223
rect 38209 12189 38243 12223
rect 40141 12189 40175 12223
rect 40325 12189 40359 12223
rect 40417 12189 40451 12223
rect 42993 12189 43027 12223
rect 43177 12189 43211 12223
rect 43272 12189 43306 12223
rect 43361 12189 43395 12223
rect 45477 12189 45511 12223
rect 46581 12189 46615 12223
rect 46765 12189 46799 12223
rect 47041 12189 47075 12223
rect 48237 12189 48271 12223
rect 48400 12189 48434 12223
rect 48500 12189 48534 12223
rect 48605 12189 48639 12223
rect 49433 12189 49467 12223
rect 49617 12189 49651 12223
rect 50537 12189 50571 12223
rect 50905 12189 50939 12223
rect 51089 12189 51123 12223
rect 52285 12189 52319 12223
rect 52469 12189 52503 12223
rect 52561 12189 52595 12223
rect 52745 12189 52779 12223
rect 53573 12189 53607 12223
rect 53941 12189 53975 12223
rect 54585 12189 54619 12223
rect 54861 12189 54895 12223
rect 55873 12189 55907 12223
rect 25237 12121 25271 12155
rect 30113 12121 30147 12155
rect 32137 12121 32171 12155
rect 33793 12121 33827 12155
rect 34989 12121 35023 12155
rect 35173 12121 35207 12155
rect 38669 12121 38703 12155
rect 45201 12121 45235 12155
rect 46673 12121 46707 12155
rect 46883 12121 46917 12155
rect 57805 12121 57839 12155
rect 24041 12053 24075 12087
rect 26617 12053 26651 12087
rect 29193 12053 29227 12087
rect 34253 12053 34287 12087
rect 35074 12053 35108 12087
rect 35725 12053 35759 12087
rect 36369 12053 36403 12087
rect 41061 12053 41095 12087
rect 41613 12053 41647 12087
rect 44189 12053 44223 12087
rect 45385 12053 45419 12087
rect 48881 12053 48915 12087
rect 50353 12053 50387 12087
rect 54769 12053 54803 12087
rect 55965 12053 55999 12087
rect 57345 12053 57379 12087
rect 24777 11849 24811 11883
rect 25513 11849 25547 11883
rect 27537 11849 27571 11883
rect 29193 11849 29227 11883
rect 31585 11849 31619 11883
rect 33517 11849 33551 11883
rect 37657 11849 37691 11883
rect 39405 11849 39439 11883
rect 40693 11849 40727 11883
rect 42073 11849 42107 11883
rect 44281 11849 44315 11883
rect 44465 11849 44499 11883
rect 45385 11849 45419 11883
rect 46857 11849 46891 11883
rect 48329 11849 48363 11883
rect 49801 11849 49835 11883
rect 50629 11849 50663 11883
rect 50813 11849 50847 11883
rect 53941 11849 53975 11883
rect 54309 11849 54343 11883
rect 55965 11849 55999 11883
rect 24133 11781 24167 11815
rect 27169 11781 27203 11815
rect 30849 11781 30883 11815
rect 31033 11781 31067 11815
rect 32413 11781 32447 11815
rect 33885 11781 33919 11815
rect 39037 11781 39071 11815
rect 39237 11781 39271 11815
rect 43729 11781 43763 11815
rect 48881 11781 48915 11815
rect 55597 11781 55631 11815
rect 55797 11781 55831 11815
rect 1869 11713 1903 11747
rect 24869 11713 24903 11747
rect 25053 11713 25087 11747
rect 25697 11713 25731 11747
rect 26065 11713 26099 11747
rect 26249 11713 26283 11747
rect 27629 11713 27663 11747
rect 28917 11713 28951 11747
rect 29285 11713 29319 11747
rect 30757 11713 30791 11747
rect 31493 11713 31527 11747
rect 31677 11713 31711 11747
rect 32321 11703 32355 11737
rect 32505 11713 32539 11747
rect 33057 11713 33091 11747
rect 33655 11713 33689 11747
rect 33793 11713 33827 11747
rect 34068 11713 34102 11747
rect 34161 11713 34195 11747
rect 34621 11713 34655 11747
rect 34713 11713 34747 11747
rect 35633 11713 35667 11747
rect 36093 11713 36127 11747
rect 36553 11713 36587 11747
rect 36737 11713 36771 11747
rect 37933 11713 37967 11747
rect 38117 11713 38151 11747
rect 40049 11713 40083 11747
rect 40233 11713 40267 11747
rect 41705 11713 41739 11747
rect 42993 11713 43027 11747
rect 43177 11713 43211 11747
rect 43453 11713 43487 11747
rect 44462 11713 44496 11747
rect 44925 11713 44959 11747
rect 45569 11713 45603 11747
rect 45753 11713 45787 11747
rect 45845 11713 45879 11747
rect 46397 11713 46431 11747
rect 46857 11713 46891 11747
rect 48605 11713 48639 11747
rect 49433 11713 49467 11747
rect 50810 11713 50844 11747
rect 51273 11713 51307 11747
rect 52009 11713 52043 11747
rect 52101 11713 52135 11747
rect 52193 11713 52227 11747
rect 52377 11713 52411 11747
rect 53849 11713 53883 11747
rect 54125 11713 54159 11747
rect 54861 11713 54895 11747
rect 55045 11713 55079 11747
rect 56977 11713 57011 11747
rect 25881 11645 25915 11679
rect 25973 11645 26007 11679
rect 27261 11645 27295 11679
rect 28733 11645 28767 11679
rect 34897 11645 34931 11679
rect 35357 11645 35391 11679
rect 35909 11645 35943 11679
rect 37841 11645 37875 11679
rect 38025 11645 38059 11679
rect 41797 11645 41831 11679
rect 44833 11645 44867 11679
rect 46673 11645 46707 11679
rect 48513 11645 48547 11679
rect 48973 11645 49007 11679
rect 49525 11645 49559 11679
rect 51181 11645 51215 11679
rect 51733 11645 51767 11679
rect 1685 11577 1719 11611
rect 2421 11577 2455 11611
rect 31033 11577 31067 11611
rect 35725 11577 35759 11611
rect 43269 11577 43303 11611
rect 45661 11577 45695 11611
rect 47777 11577 47811 11611
rect 54861 11577 54895 11611
rect 24593 11509 24627 11543
rect 27353 11509 27387 11543
rect 28089 11509 28123 11543
rect 29837 11509 29871 11543
rect 34805 11509 34839 11543
rect 35817 11509 35851 11543
rect 36737 11509 36771 11543
rect 39221 11509 39255 11543
rect 40233 11509 40267 11543
rect 43361 11509 43395 11543
rect 46535 11509 46569 11543
rect 49433 11509 49467 11543
rect 52929 11509 52963 11543
rect 55781 11509 55815 11543
rect 56517 11509 56551 11543
rect 58173 11509 58207 11543
rect 24961 11305 24995 11339
rect 25605 11305 25639 11339
rect 27445 11305 27479 11339
rect 28273 11305 28307 11339
rect 29837 11305 29871 11339
rect 30573 11305 30607 11339
rect 32137 11305 32171 11339
rect 32965 11305 32999 11339
rect 33885 11305 33919 11339
rect 34345 11305 34379 11339
rect 36093 11305 36127 11339
rect 37749 11305 37783 11339
rect 38669 11305 38703 11339
rect 40785 11305 40819 11339
rect 42349 11305 42383 11339
rect 43085 11305 43119 11339
rect 44005 11305 44039 11339
rect 46397 11305 46431 11339
rect 48329 11305 48363 11339
rect 49617 11305 49651 11339
rect 50997 11305 51031 11339
rect 53021 11305 53055 11339
rect 54401 11305 54435 11339
rect 55873 11305 55907 11339
rect 58081 11305 58115 11339
rect 26341 11237 26375 11271
rect 36553 11237 36587 11271
rect 41245 11237 41279 11271
rect 51733 11237 51767 11271
rect 52837 11237 52871 11271
rect 24593 11169 24627 11203
rect 30849 11169 30883 11203
rect 40141 11169 40175 11203
rect 45293 11169 45327 11203
rect 47409 11169 47443 11203
rect 47501 11169 47535 11203
rect 48973 11169 49007 11203
rect 52101 11169 52135 11203
rect 53941 11169 53975 11203
rect 54217 11169 54251 11203
rect 24777 11101 24811 11135
rect 25421 11101 25455 11135
rect 25605 11101 25639 11135
rect 27813 11101 27847 11135
rect 28457 11101 28491 11135
rect 28641 11101 28675 11135
rect 28733 11101 28767 11135
rect 29745 11101 29779 11135
rect 29929 11101 29963 11135
rect 30757 11101 30791 11135
rect 30941 11101 30975 11135
rect 31069 11101 31103 11135
rect 32045 11101 32079 11135
rect 32229 11101 32263 11135
rect 32689 11079 32723 11113
rect 33793 11101 33827 11135
rect 34161 11101 34195 11135
rect 35541 11101 35575 11135
rect 36829 11101 36863 11135
rect 37289 11101 37323 11135
rect 37565 11101 37599 11135
rect 38853 11101 38887 11135
rect 40417 11101 40451 11135
rect 42901 11101 42935 11135
rect 43085 11101 43119 11135
rect 43545 11101 43579 11135
rect 43821 11101 43855 11135
rect 45193 11101 45227 11135
rect 47317 11101 47351 11135
rect 47593 11101 47627 11135
rect 48329 11101 48363 11135
rect 48513 11101 48547 11135
rect 50353 11101 50387 11135
rect 50537 11101 50571 11135
rect 50629 11101 50663 11135
rect 50721 11101 50755 11135
rect 51917 11101 51951 11135
rect 52009 11101 52043 11135
rect 52193 11101 52227 11135
rect 52377 11101 52411 11135
rect 54033 11101 54067 11135
rect 54125 11101 54159 11135
rect 55505 11101 55539 11135
rect 56333 11101 56367 11135
rect 56517 11101 56551 11135
rect 27629 11033 27663 11067
rect 32781 11033 32815 11067
rect 32965 11033 32999 11067
rect 36553 11033 36587 11067
rect 36737 11033 36771 11067
rect 39313 11033 39347 11067
rect 40325 11033 40359 11067
rect 43637 11033 43671 11067
rect 44557 11033 44591 11067
rect 53205 11033 53239 11067
rect 54861 11033 54895 11067
rect 55689 11033 55723 11067
rect 56425 11033 56459 11067
rect 26893 10965 26927 10999
rect 34897 10965 34931 10999
rect 37381 10965 37415 10999
rect 41797 10965 41831 10999
rect 45845 10965 45879 10999
rect 47777 10965 47811 10999
rect 53005 10965 53039 10999
rect 56977 10965 57011 10999
rect 57529 10965 57563 10999
rect 28733 10761 28767 10795
rect 30297 10761 30331 10795
rect 31033 10761 31067 10795
rect 32321 10761 32355 10795
rect 33885 10761 33919 10795
rect 35081 10761 35115 10795
rect 38209 10761 38243 10795
rect 39313 10761 39347 10795
rect 49433 10761 49467 10795
rect 50537 10761 50571 10795
rect 52193 10761 52227 10795
rect 54033 10761 54067 10795
rect 55045 10761 55079 10795
rect 57437 10761 57471 10795
rect 24225 10693 24259 10727
rect 28641 10693 28675 10727
rect 31201 10693 31235 10727
rect 31401 10693 31435 10727
rect 42809 10693 42843 10727
rect 48053 10693 48087 10727
rect 48697 10693 48731 10727
rect 53021 10693 53055 10727
rect 24961 10625 24995 10659
rect 26249 10625 26283 10659
rect 27353 10625 27387 10659
rect 27629 10625 27663 10659
rect 29837 10625 29871 10659
rect 29929 10625 29963 10659
rect 30093 10625 30127 10659
rect 32597 10625 32631 10659
rect 34161 10625 34195 10659
rect 35449 10625 35483 10659
rect 35541 10625 35575 10659
rect 36553 10625 36587 10659
rect 36921 10625 36955 10659
rect 37565 10625 37599 10659
rect 37749 10625 37783 10659
rect 38577 10625 38611 10659
rect 39221 10625 39255 10659
rect 39405 10625 39439 10659
rect 40693 10625 40727 10659
rect 41245 10625 41279 10659
rect 44281 10625 44315 10659
rect 45293 10625 45327 10659
rect 45477 10625 45511 10659
rect 46121 10625 46155 10659
rect 46489 10625 46523 10659
rect 46949 10625 46983 10659
rect 47777 10625 47811 10659
rect 47869 10625 47903 10659
rect 48605 10625 48639 10659
rect 48881 10625 48915 10659
rect 49801 10625 49835 10659
rect 50261 10625 50295 10659
rect 50353 10625 50387 10659
rect 51641 10625 51675 10659
rect 52101 10625 52135 10659
rect 52285 10625 52319 10659
rect 52929 10625 52963 10659
rect 53113 10625 53147 10659
rect 54217 10625 54251 10659
rect 54309 10625 54343 10659
rect 54585 10625 54619 10659
rect 56241 10625 56275 10659
rect 24685 10557 24719 10591
rect 27445 10557 27479 10591
rect 28825 10557 28859 10591
rect 32505 10557 32539 10591
rect 32689 10557 32723 10591
rect 32781 10557 32815 10591
rect 34069 10557 34103 10591
rect 34253 10557 34287 10591
rect 34345 10557 34379 10591
rect 35265 10557 35299 10591
rect 35357 10557 35391 10591
rect 37657 10557 37691 10591
rect 38393 10557 38427 10591
rect 38485 10557 38519 10591
rect 38669 10557 38703 10591
rect 44465 10557 44499 10591
rect 46213 10557 46247 10591
rect 46765 10557 46799 10591
rect 49709 10557 49743 10591
rect 50537 10557 50571 10591
rect 51549 10557 51583 10591
rect 54493 10557 54527 10591
rect 24777 10489 24811 10523
rect 27537 10489 27571 10523
rect 36369 10489 36403 10523
rect 46489 10489 46523 10523
rect 47777 10489 47811 10523
rect 48881 10489 48915 10523
rect 55965 10489 55999 10523
rect 24869 10421 24903 10455
rect 25697 10421 25731 10455
rect 26433 10421 26467 10455
rect 27169 10421 27203 10455
rect 28273 10421 28307 10455
rect 31226 10421 31260 10455
rect 33425 10421 33459 10455
rect 36737 10421 36771 10455
rect 43269 10421 43303 10455
rect 44097 10421 44131 10455
rect 45385 10421 45419 10455
rect 49801 10421 49835 10455
rect 51273 10421 51307 10455
rect 51457 10421 51491 10455
rect 56793 10421 56827 10455
rect 58081 10421 58115 10455
rect 24593 10217 24627 10251
rect 26249 10217 26283 10251
rect 26801 10217 26835 10251
rect 28457 10217 28491 10251
rect 29193 10217 29227 10251
rect 29929 10217 29963 10251
rect 30573 10217 30607 10251
rect 31585 10217 31619 10251
rect 38301 10217 38335 10251
rect 38485 10217 38519 10251
rect 38945 10217 38979 10251
rect 43177 10217 43211 10251
rect 43821 10217 43855 10251
rect 44005 10217 44039 10251
rect 45937 10217 45971 10251
rect 47225 10217 47259 10251
rect 47685 10217 47719 10251
rect 49157 10217 49191 10251
rect 50813 10217 50847 10251
rect 52377 10217 52411 10251
rect 53205 10217 53239 10251
rect 53849 10217 53883 10251
rect 54493 10217 54527 10251
rect 36829 10149 36863 10183
rect 41613 10149 41647 10183
rect 42625 10149 42659 10183
rect 45385 10149 45419 10183
rect 47961 10149 47995 10183
rect 51457 10149 51491 10183
rect 51549 10149 51583 10183
rect 58173 10149 58207 10183
rect 32505 10081 32539 10115
rect 33885 10081 33919 10115
rect 36553 10081 36587 10115
rect 42165 10081 42199 10115
rect 43361 10081 43395 10115
rect 45293 10081 45327 10115
rect 48053 10081 48087 10115
rect 49341 10081 49375 10115
rect 23857 10013 23891 10047
rect 24041 10013 24075 10047
rect 24869 10013 24903 10047
rect 25329 10013 25363 10047
rect 25513 10013 25547 10047
rect 25789 10013 25823 10047
rect 26430 10013 26464 10047
rect 26893 10013 26927 10047
rect 27813 10013 27847 10047
rect 27997 10013 28031 10047
rect 28089 10013 28123 10047
rect 28227 10013 28261 10047
rect 29745 10013 29779 10047
rect 29929 10013 29963 10047
rect 30389 10013 30423 10047
rect 30573 10013 30607 10047
rect 31493 10013 31527 10047
rect 31677 10013 31711 10047
rect 32413 10013 32447 10047
rect 32597 10013 32631 10047
rect 33057 10013 33091 10047
rect 33253 10013 33287 10047
rect 33793 10013 33827 10047
rect 34069 10013 34103 10047
rect 34161 10013 34195 10047
rect 35357 10013 35391 10047
rect 35817 10013 35851 10047
rect 36369 10013 36403 10047
rect 36921 10013 36955 10047
rect 39129 10013 39163 10047
rect 39221 10013 39255 10047
rect 40049 10013 40083 10047
rect 40233 10013 40267 10047
rect 41337 10013 41371 10047
rect 42257 10013 42291 10047
rect 43085 10013 43119 10047
rect 45756 10013 45790 10047
rect 46857 10013 46891 10047
rect 47041 10013 47075 10047
rect 47869 10013 47903 10047
rect 48145 10013 48179 10047
rect 48329 10013 48363 10047
rect 49433 10013 49467 10047
rect 50629 10013 50663 10047
rect 50813 10013 50847 10047
rect 51365 10013 51399 10047
rect 51641 10013 51675 10047
rect 53113 10013 53147 10047
rect 53297 10013 53331 10047
rect 53757 10013 53791 10047
rect 53941 10013 53975 10047
rect 56149 10013 56183 10047
rect 56425 10013 56459 10047
rect 24593 9945 24627 9979
rect 24777 9945 24811 9979
rect 33149 9945 33183 9979
rect 33701 9945 33735 9979
rect 38117 9945 38151 9979
rect 38317 9945 38351 9979
rect 40417 9945 40451 9979
rect 41613 9945 41647 9979
rect 43361 9945 43395 9979
rect 43989 9945 44023 9979
rect 44189 9945 44223 9979
rect 49709 9945 49743 9979
rect 49801 9945 49835 9979
rect 51825 9945 51859 9979
rect 24041 9877 24075 9911
rect 25697 9877 25731 9911
rect 26433 9877 26467 9911
rect 41429 9877 41463 9911
rect 45753 9877 45787 9911
rect 55965 9877 55999 9911
rect 57069 9877 57103 9911
rect 57621 9877 57655 9911
rect 27445 9673 27479 9707
rect 34161 9673 34195 9707
rect 36369 9673 36403 9707
rect 39773 9673 39807 9707
rect 56333 9673 56367 9707
rect 23765 9605 23799 9639
rect 24869 9605 24903 9639
rect 27353 9605 27387 9639
rect 28457 9605 28491 9639
rect 30757 9605 30791 9639
rect 32781 9605 32815 9639
rect 36001 9605 36035 9639
rect 36201 9605 36235 9639
rect 40877 9605 40911 9639
rect 44373 9605 44407 9639
rect 44557 9605 44591 9639
rect 45661 9605 45695 9639
rect 48697 9605 48731 9639
rect 50261 9605 50295 9639
rect 51917 9605 51951 9639
rect 53113 9605 53147 9639
rect 53205 9605 53239 9639
rect 55781 9605 55815 9639
rect 58081 9605 58115 9639
rect 28641 9537 28675 9571
rect 28733 9537 28767 9571
rect 28917 9537 28951 9571
rect 29019 9527 29053 9561
rect 29653 9537 29687 9571
rect 29837 9537 29871 9571
rect 30113 9537 30147 9571
rect 30941 9537 30975 9571
rect 31033 9537 31067 9571
rect 31217 9537 31251 9571
rect 31309 9537 31343 9571
rect 32948 9537 32982 9571
rect 33057 9537 33091 9571
rect 33333 9537 33367 9571
rect 33793 9537 33827 9571
rect 33977 9537 34011 9571
rect 34897 9537 34931 9571
rect 35081 9537 35115 9571
rect 37473 9537 37507 9571
rect 38209 9537 38243 9571
rect 39589 9537 39623 9571
rect 43637 9537 43671 9571
rect 44097 9537 44131 9571
rect 45109 9537 45143 9571
rect 45845 9537 45879 9571
rect 46029 9537 46063 9571
rect 46121 9537 46155 9571
rect 48145 9537 48179 9571
rect 48911 9537 48945 9571
rect 49157 9537 49191 9571
rect 52101 9537 52135 9571
rect 53021 9537 53055 9571
rect 53389 9537 53423 9571
rect 53481 9537 53515 9571
rect 54217 9537 54251 9571
rect 54459 9537 54493 9571
rect 56425 9537 56459 9571
rect 24317 9469 24351 9503
rect 26065 9469 26099 9503
rect 27721 9469 27755 9503
rect 29929 9469 29963 9503
rect 36829 9469 36863 9503
rect 37749 9469 37783 9503
rect 43545 9469 43579 9503
rect 45753 9469 45787 9503
rect 52377 9469 52411 9503
rect 52929 9469 52963 9503
rect 54769 9469 54803 9503
rect 54861 9469 54895 9503
rect 27537 9401 27571 9435
rect 29469 9401 29503 9435
rect 29745 9401 29779 9435
rect 33241 9401 33275 9435
rect 38945 9401 38979 9435
rect 40325 9401 40359 9435
rect 41521 9401 41555 9435
rect 41981 9401 42015 9435
rect 43269 9401 43303 9435
rect 47961 9401 47995 9435
rect 49065 9401 49099 9435
rect 49709 9401 49743 9435
rect 52285 9401 52319 9435
rect 55321 9401 55355 9435
rect 55505 9401 55539 9435
rect 56885 9401 56919 9435
rect 24961 9333 24995 9367
rect 26617 9333 26651 9367
rect 27629 9333 27663 9367
rect 34897 9333 34931 9367
rect 35265 9333 35299 9367
rect 36185 9333 36219 9367
rect 37565 9333 37599 9367
rect 37657 9333 37691 9367
rect 38393 9333 38427 9367
rect 42625 9333 42659 9367
rect 43637 9333 43671 9367
rect 44346 9333 44380 9367
rect 46673 9333 46707 9367
rect 47225 9333 47259 9367
rect 50721 9333 50755 9367
rect 51365 9333 51399 9367
rect 57437 9333 57471 9367
rect 26157 9129 26191 9163
rect 30389 9129 30423 9163
rect 30757 9129 30791 9163
rect 32413 9129 32447 9163
rect 32965 9129 32999 9163
rect 33425 9129 33459 9163
rect 33793 9129 33827 9163
rect 35633 9129 35667 9163
rect 37289 9129 37323 9163
rect 38669 9129 38703 9163
rect 38853 9129 38887 9163
rect 39405 9129 39439 9163
rect 45661 9129 45695 9163
rect 49157 9129 49191 9163
rect 50813 9129 50847 9163
rect 53205 9129 53239 9163
rect 55597 9129 55631 9163
rect 56149 9129 56183 9163
rect 26065 9061 26099 9095
rect 27537 9061 27571 9095
rect 29009 9061 29043 9095
rect 29929 9061 29963 9095
rect 31493 9061 31527 9095
rect 37749 9061 37783 9095
rect 41245 9061 41279 9095
rect 42441 9061 42475 9095
rect 47041 9061 47075 9095
rect 50905 9061 50939 9095
rect 51733 9061 51767 9095
rect 54861 9061 54895 9095
rect 58265 9061 58299 9095
rect 24685 8993 24719 9027
rect 25237 8993 25271 9027
rect 27997 8993 28031 9027
rect 30481 8993 30515 9027
rect 32689 8993 32723 9027
rect 36829 8993 36863 9027
rect 41337 8993 41371 9027
rect 53941 8993 53975 9027
rect 54033 8993 54067 9027
rect 25973 8925 26007 8959
rect 26249 8925 26283 8959
rect 26433 8925 26467 8959
rect 27721 8925 27755 8959
rect 27905 8925 27939 8959
rect 28089 8925 28123 8959
rect 28273 8925 28307 8959
rect 29193 8925 29227 8959
rect 29745 8925 29779 8959
rect 29929 8925 29963 8959
rect 30389 8925 30423 8959
rect 31493 8925 31527 8959
rect 31677 8925 31711 8959
rect 32781 8925 32815 8959
rect 33425 8925 33459 8959
rect 33609 8925 33643 8959
rect 34897 8925 34931 8959
rect 35081 8925 35115 8959
rect 35725 8925 35759 8959
rect 36921 8925 36955 8959
rect 37105 8925 37139 8959
rect 38485 8925 38519 8959
rect 38761 8925 38795 8959
rect 40233 8925 40267 8959
rect 40601 8925 40635 8959
rect 41061 8925 41095 8959
rect 41153 8925 41187 8959
rect 42073 8925 42107 8959
rect 42166 8925 42200 8959
rect 45845 8925 45879 8959
rect 46121 8925 46155 8959
rect 46305 8925 46339 8959
rect 46765 8925 46799 8959
rect 47685 8925 47719 8959
rect 48605 8925 48639 8959
rect 51917 8925 51951 8959
rect 53021 8925 53055 8959
rect 53205 8925 53239 8959
rect 53665 8925 53699 8959
rect 53849 8925 53883 8959
rect 54125 8925 54159 8959
rect 54309 8925 54343 8959
rect 57161 8925 57195 8959
rect 32321 8857 32355 8891
rect 36277 8857 36311 8891
rect 38393 8857 38427 8891
rect 40325 8857 40359 8891
rect 40417 8857 40451 8891
rect 42993 8857 43027 8891
rect 44189 8857 44223 8891
rect 44557 8857 44591 8891
rect 45937 8857 45971 8891
rect 46029 8857 46063 8891
rect 46857 8857 46891 8891
rect 47041 8857 47075 8891
rect 48237 8857 48271 8891
rect 51273 8857 51307 8891
rect 52101 8857 52135 8891
rect 24041 8789 24075 8823
rect 25697 8789 25731 8823
rect 26985 8789 27019 8823
rect 34345 8789 34379 8823
rect 34989 8789 35023 8823
rect 40049 8789 40083 8823
rect 43545 8789 43579 8823
rect 47593 8789 47627 8823
rect 49709 8789 49743 8823
rect 56701 8789 56735 8823
rect 57713 8789 57747 8823
rect 25053 8585 25087 8619
rect 27813 8585 27847 8619
rect 28733 8585 28767 8619
rect 32689 8585 32723 8619
rect 37565 8585 37599 8619
rect 38945 8585 38979 8619
rect 44005 8585 44039 8619
rect 47869 8585 47903 8619
rect 48789 8585 48823 8619
rect 50721 8585 50755 8619
rect 54677 8585 54711 8619
rect 58081 8585 58115 8619
rect 25605 8517 25639 8551
rect 25697 8517 25731 8551
rect 26617 8517 26651 8551
rect 29837 8517 29871 8551
rect 30757 8517 30791 8551
rect 45661 8517 45695 8551
rect 46213 8517 46247 8551
rect 51641 8517 51675 8551
rect 56977 8517 57011 8551
rect 25329 8449 25363 8483
rect 27169 8449 27203 8483
rect 27625 8449 27659 8483
rect 28917 8449 28951 8483
rect 29193 8449 29227 8483
rect 29745 8449 29779 8483
rect 29929 8449 29963 8483
rect 30573 8449 30607 8483
rect 30941 8449 30975 8483
rect 31217 8449 31251 8483
rect 31769 8449 31803 8483
rect 32689 8449 32723 8483
rect 33865 8449 33899 8483
rect 33977 8449 34011 8483
rect 34074 8449 34108 8483
rect 34253 8449 34287 8483
rect 35173 8449 35207 8483
rect 35265 8449 35299 8483
rect 35449 8449 35483 8483
rect 35633 8449 35667 8483
rect 36369 8449 36403 8483
rect 36461 8449 36495 8483
rect 36553 8449 36587 8483
rect 36737 8449 36771 8483
rect 37749 8449 37783 8483
rect 37933 8449 37967 8483
rect 38761 8449 38795 8483
rect 39405 8449 39439 8483
rect 39589 8449 39623 8483
rect 40601 8449 40635 8483
rect 41429 8449 41463 8483
rect 41797 8449 41831 8483
rect 42073 8449 42107 8483
rect 42717 8449 42751 8483
rect 43545 8449 43579 8483
rect 44373 8449 44407 8483
rect 45201 8449 45235 8483
rect 45477 8449 45511 8483
rect 46121 8449 46155 8483
rect 46305 8449 46339 8483
rect 46949 8449 46983 8483
rect 47133 8449 47167 8483
rect 48053 8449 48087 8483
rect 49617 8449 49651 8483
rect 49709 8449 49743 8483
rect 50077 8449 50111 8483
rect 51825 8449 51859 8483
rect 52009 8449 52043 8483
rect 52101 8449 52135 8483
rect 52929 8449 52963 8483
rect 53389 8449 53423 8483
rect 54677 8449 54711 8483
rect 55321 8449 55355 8483
rect 55413 8449 55447 8483
rect 55781 8449 55815 8483
rect 56425 8449 56459 8483
rect 23949 8381 23983 8415
rect 24501 8381 24535 8415
rect 25217 8381 25251 8415
rect 27353 8381 27387 8415
rect 27445 8381 27479 8415
rect 29009 8381 29043 8415
rect 30389 8381 30423 8415
rect 32321 8381 32355 8415
rect 32873 8381 32907 8415
rect 34989 8381 35023 8415
rect 38485 8381 38519 8415
rect 40325 8381 40359 8415
rect 43177 8381 43211 8415
rect 44465 8381 44499 8415
rect 44557 8381 44591 8415
rect 48329 8381 48363 8415
rect 49801 8381 49835 8415
rect 49893 8381 49927 8415
rect 50537 8381 50571 8415
rect 50905 8381 50939 8415
rect 53665 8381 53699 8415
rect 27537 8313 27571 8347
rect 29101 8313 29135 8347
rect 35357 8313 35391 8347
rect 39773 8313 39807 8347
rect 40785 8313 40819 8347
rect 41521 8313 41555 8347
rect 47133 8313 47167 8347
rect 48237 8313 48271 8347
rect 49433 8313 49467 8347
rect 54217 8313 54251 8347
rect 55413 8313 55447 8347
rect 33609 8245 33643 8279
rect 36093 8245 36127 8279
rect 38577 8245 38611 8279
rect 40417 8245 40451 8279
rect 45293 8245 45327 8279
rect 50905 8245 50939 8279
rect 24593 8041 24627 8075
rect 27445 8041 27479 8075
rect 29929 8041 29963 8075
rect 33241 8041 33275 8075
rect 35265 8041 35299 8075
rect 35817 8041 35851 8075
rect 36001 8041 36035 8075
rect 36829 8041 36863 8075
rect 38761 8041 38795 8075
rect 40417 8041 40451 8075
rect 40969 8041 41003 8075
rect 42073 8041 42107 8075
rect 45845 8041 45879 8075
rect 48329 8041 48363 8075
rect 49801 8041 49835 8075
rect 51825 8041 51859 8075
rect 52653 8041 52687 8075
rect 56149 8041 56183 8075
rect 57437 8041 57471 8075
rect 25789 7973 25823 8007
rect 27077 7973 27111 8007
rect 33793 7973 33827 8007
rect 38945 7973 38979 8007
rect 42809 7973 42843 8007
rect 53573 7973 53607 8007
rect 55873 7973 55907 8007
rect 55965 7973 55999 8007
rect 25513 7905 25547 7939
rect 35173 7905 35207 7939
rect 35357 7905 35391 7939
rect 39221 7905 39255 7939
rect 49433 7905 49467 7939
rect 50721 7905 50755 7939
rect 56057 7905 56091 7939
rect 25237 7837 25271 7871
rect 25396 7837 25430 7871
rect 26249 7837 26283 7871
rect 26433 7837 26467 7871
rect 26985 7837 27019 7871
rect 27261 7837 27295 7871
rect 27997 7837 28031 7871
rect 28549 7837 28583 7871
rect 28825 7837 28859 7871
rect 29745 7837 29779 7871
rect 29837 7837 29871 7871
rect 31401 7837 31435 7871
rect 31769 7837 31803 7871
rect 32137 7837 32171 7871
rect 33149 7837 33183 7871
rect 33241 7837 33275 7871
rect 33793 7837 33827 7871
rect 34069 7837 34103 7871
rect 35081 7837 35115 7871
rect 36001 7837 36035 7871
rect 36185 7837 36219 7871
rect 36737 7837 36771 7871
rect 37749 7837 37783 7871
rect 38025 7837 38059 7871
rect 40141 7837 40175 7871
rect 42625 7837 42659 7871
rect 42809 7837 42843 7871
rect 46581 7837 46615 7871
rect 46673 7837 46707 7871
rect 46869 7837 46903 7871
rect 46959 7837 46993 7871
rect 47685 7837 47719 7871
rect 47869 7837 47903 7871
rect 47961 7837 47995 7871
rect 48053 7837 48087 7871
rect 49341 7837 49375 7871
rect 49525 7837 49559 7871
rect 49617 7837 49651 7871
rect 51273 7837 51307 7871
rect 51365 7837 51399 7871
rect 51549 7837 51583 7871
rect 51641 7837 51675 7871
rect 52837 7837 52871 7871
rect 53021 7837 53055 7871
rect 53113 7837 53147 7871
rect 53757 7837 53791 7871
rect 53941 7837 53975 7871
rect 54401 7837 54435 7871
rect 54585 7837 54619 7871
rect 55505 7837 55539 7871
rect 28457 7769 28491 7803
rect 43821 7769 43855 7803
rect 50445 7769 50479 7803
rect 30113 7701 30147 7735
rect 30665 7701 30699 7735
rect 31309 7701 31343 7735
rect 33977 7701 34011 7735
rect 38209 7701 38243 7735
rect 41521 7701 41555 7735
rect 43913 7701 43947 7735
rect 45293 7701 45327 7735
rect 46397 7701 46431 7735
rect 54493 7701 54527 7735
rect 56885 7701 56919 7735
rect 57989 7701 58023 7735
rect 24777 7497 24811 7531
rect 25789 7497 25823 7531
rect 27169 7497 27203 7531
rect 30297 7497 30331 7531
rect 31401 7497 31435 7531
rect 34529 7497 34563 7531
rect 35633 7497 35667 7531
rect 36829 7497 36863 7531
rect 38393 7497 38427 7531
rect 40785 7497 40819 7531
rect 44205 7497 44239 7531
rect 44833 7497 44867 7531
rect 46029 7497 46063 7531
rect 51365 7497 51399 7531
rect 53021 7497 53055 7531
rect 54217 7497 54251 7531
rect 56609 7497 56643 7531
rect 33057 7429 33091 7463
rect 37473 7429 37507 7463
rect 39497 7429 39531 7463
rect 44005 7429 44039 7463
rect 46305 7429 46339 7463
rect 46397 7429 46431 7463
rect 47133 7429 47167 7463
rect 51917 7429 51951 7463
rect 52285 7429 52319 7463
rect 24685 7361 24719 7395
rect 24961 7361 24995 7395
rect 25973 7361 26007 7395
rect 26065 7361 26099 7395
rect 26249 7361 26283 7395
rect 26341 7361 26375 7395
rect 27353 7361 27387 7395
rect 27629 7361 27663 7395
rect 27813 7361 27847 7395
rect 28641 7361 28675 7395
rect 29469 7361 29503 7395
rect 29653 7361 29687 7395
rect 30481 7361 30515 7395
rect 30665 7361 30699 7395
rect 31585 7361 31619 7395
rect 33701 7361 33735 7395
rect 33793 7361 33827 7395
rect 33977 7361 34011 7395
rect 36461 7361 36495 7395
rect 36645 7361 36679 7395
rect 38209 7361 38243 7395
rect 38301 7361 38335 7395
rect 39129 7361 39163 7395
rect 40141 7361 40175 7395
rect 40969 7361 41003 7395
rect 42901 7361 42935 7395
rect 42993 7361 43027 7395
rect 45293 7361 45327 7395
rect 46213 7361 46247 7395
rect 46535 7361 46569 7395
rect 47961 7361 47995 7395
rect 48145 7361 48179 7395
rect 48789 7361 48823 7395
rect 49709 7361 49743 7395
rect 49801 7361 49835 7395
rect 50997 7361 51031 7395
rect 51457 7361 51491 7395
rect 52929 7361 52963 7395
rect 53205 7361 53239 7395
rect 54493 7361 54527 7395
rect 54677 7361 54711 7395
rect 54861 7361 54895 7395
rect 58081 7361 58115 7395
rect 27537 7293 27571 7327
rect 28365 7293 28399 7327
rect 29009 7293 29043 7327
rect 30573 7293 30607 7327
rect 30757 7293 30791 7327
rect 32505 7293 32539 7327
rect 32689 7293 32723 7327
rect 35173 7293 35207 7327
rect 38025 7293 38059 7327
rect 38577 7293 38611 7327
rect 40325 7293 40359 7327
rect 41153 7293 41187 7327
rect 42809 7293 42843 7327
rect 43085 7293 43119 7327
rect 46673 7293 46707 7327
rect 47777 7293 47811 7327
rect 48237 7293 48271 7327
rect 49617 7293 49651 7327
rect 49893 7293 49927 7327
rect 51089 7293 51123 7327
rect 54585 7293 54619 7327
rect 27445 7225 27479 7259
rect 32919 7225 32953 7259
rect 33885 7225 33919 7259
rect 35541 7225 35575 7259
rect 39957 7225 39991 7259
rect 41613 7225 41647 7259
rect 48881 7225 48915 7259
rect 51181 7225 51215 7259
rect 24961 7157 24995 7191
rect 32781 7157 32815 7191
rect 33517 7157 33551 7191
rect 42625 7157 42659 7191
rect 44189 7157 44223 7191
rect 44373 7157 44407 7191
rect 45201 7157 45235 7191
rect 49433 7157 49467 7191
rect 50721 7157 50755 7191
rect 53389 7157 53423 7191
rect 54769 7157 54803 7191
rect 55505 7157 55539 7191
rect 55965 7157 55999 7191
rect 57069 7157 57103 7191
rect 58265 7157 58299 7191
rect 26801 6953 26835 6987
rect 28089 6953 28123 6987
rect 33793 6953 33827 6987
rect 34989 6953 35023 6987
rect 41889 6953 41923 6987
rect 43821 6953 43855 6987
rect 47225 6953 47259 6987
rect 48145 6953 48179 6987
rect 48513 6953 48547 6987
rect 49525 6953 49559 6987
rect 56333 6953 56367 6987
rect 58081 6953 58115 6987
rect 35081 6885 35115 6919
rect 41337 6885 41371 6919
rect 46489 6885 46523 6919
rect 50445 6885 50479 6919
rect 54677 6885 54711 6919
rect 28273 6817 28307 6851
rect 29837 6817 29871 6851
rect 30297 6817 30331 6851
rect 30665 6817 30699 6851
rect 33057 6817 33091 6851
rect 33149 6817 33183 6851
rect 34161 6817 34195 6851
rect 35449 6817 35483 6851
rect 37105 6817 37139 6851
rect 42533 6817 42567 6851
rect 42993 6817 43027 6851
rect 47409 6817 47443 6851
rect 49065 6817 49099 6851
rect 51825 6817 51859 6851
rect 55505 6817 55539 6851
rect 56885 6817 56919 6851
rect 57437 6817 57471 6851
rect 24041 6749 24075 6783
rect 25053 6749 25087 6783
rect 25146 6749 25180 6783
rect 25329 6749 25363 6783
rect 25559 6749 25593 6783
rect 26525 6749 26559 6783
rect 27353 6749 27387 6783
rect 27537 6749 27571 6783
rect 28365 6749 28399 6783
rect 29193 6749 29227 6783
rect 30481 6749 30515 6783
rect 30757 6749 30791 6783
rect 30849 6749 30883 6783
rect 31033 6749 31067 6783
rect 31493 6749 31527 6783
rect 31861 6749 31895 6783
rect 31953 6749 31987 6783
rect 32690 6749 32724 6783
rect 32781 6749 32815 6783
rect 33977 6749 34011 6783
rect 36093 6749 36127 6783
rect 36277 6749 36311 6783
rect 37565 6749 37599 6783
rect 38025 6749 38059 6783
rect 39497 6749 39531 6783
rect 40233 6749 40267 6783
rect 41153 6749 41187 6783
rect 41429 6749 41463 6783
rect 42625 6749 42659 6783
rect 44465 6749 44499 6783
rect 45477 6749 45511 6783
rect 45845 6749 45879 6783
rect 47317 6749 47351 6783
rect 47593 6749 47627 6783
rect 47685 6749 47719 6783
rect 48605 6749 48639 6783
rect 49249 6749 49283 6783
rect 49341 6749 49375 6783
rect 49617 6749 49651 6783
rect 50353 6749 50387 6783
rect 50621 6749 50655 6783
rect 51733 6749 51767 6783
rect 51917 6749 51951 6783
rect 52561 6749 52595 6783
rect 55689 6749 55723 6783
rect 55781 6749 55815 6783
rect 58265 6749 58299 6783
rect 25421 6681 25455 6715
rect 26617 6681 26651 6715
rect 26801 6681 26835 6715
rect 27261 6681 27295 6715
rect 28089 6681 28123 6715
rect 40969 6681 41003 6715
rect 43913 6681 43947 6715
rect 45661 6681 45695 6715
rect 45753 6681 45787 6715
rect 52377 6681 52411 6715
rect 53297 6681 53331 6715
rect 54861 6681 54895 6715
rect 25697 6613 25731 6647
rect 28549 6613 28583 6647
rect 31769 6613 31803 6647
rect 32505 6613 32539 6647
rect 36277 6613 36311 6647
rect 39313 6613 39347 6647
rect 40417 6613 40451 6647
rect 46029 6613 46063 6647
rect 50813 6613 50847 6647
rect 52745 6613 52779 6647
rect 53389 6613 53423 6647
rect 24133 6409 24167 6443
rect 27169 6409 27203 6443
rect 29009 6409 29043 6443
rect 29653 6409 29687 6443
rect 31033 6409 31067 6443
rect 31769 6409 31803 6443
rect 32505 6409 32539 6443
rect 33885 6409 33919 6443
rect 40509 6409 40543 6443
rect 41153 6409 41187 6443
rect 43913 6409 43947 6443
rect 46121 6409 46155 6443
rect 49893 6409 49927 6443
rect 55045 6409 55079 6443
rect 58173 6409 58207 6443
rect 25605 6341 25639 6375
rect 30297 6341 30331 6375
rect 30481 6341 30515 6375
rect 33241 6341 33275 6375
rect 36461 6341 36495 6375
rect 38857 6341 38891 6375
rect 45385 6341 45419 6375
rect 52193 6341 52227 6375
rect 52377 6341 52411 6375
rect 54953 6341 54987 6375
rect 57529 6341 57563 6375
rect 24593 6273 24627 6307
rect 25329 6273 25363 6307
rect 25881 6273 25915 6307
rect 26065 6273 26099 6307
rect 28733 6273 28767 6307
rect 30113 6273 30147 6307
rect 30941 6273 30975 6307
rect 31125 6273 31159 6307
rect 32321 6273 32355 6307
rect 33701 6273 33735 6307
rect 34069 6273 34103 6307
rect 34345 6273 34379 6307
rect 35081 6273 35115 6307
rect 36277 6273 36311 6307
rect 36921 6273 36955 6307
rect 37565 6273 37599 6307
rect 38761 6273 38795 6307
rect 38945 6273 38979 6307
rect 39129 6273 39163 6307
rect 39865 6273 39899 6307
rect 40417 6273 40451 6307
rect 40601 6273 40635 6307
rect 42625 6273 42659 6307
rect 45661 6273 45695 6307
rect 46305 6273 46339 6307
rect 46581 6273 46615 6307
rect 46765 6273 46799 6307
rect 48053 6273 48087 6307
rect 48513 6273 48547 6307
rect 49433 6273 49467 6307
rect 50077 6273 50111 6307
rect 50169 6273 50203 6307
rect 50353 6273 50387 6307
rect 50537 6273 50571 6307
rect 51181 6273 51215 6307
rect 51273 6273 51307 6307
rect 53113 6273 53147 6307
rect 53389 6273 53423 6307
rect 54125 6273 54159 6307
rect 24869 6205 24903 6239
rect 26617 6205 26651 6239
rect 35265 6205 35299 6239
rect 37841 6205 37875 6239
rect 42901 6205 42935 6239
rect 50261 6205 50295 6239
rect 50997 6205 51031 6239
rect 52929 6205 52963 6239
rect 38577 6137 38611 6171
rect 41613 6137 41647 6171
rect 48789 6137 48823 6171
rect 52009 6137 52043 6171
rect 54309 6137 54343 6171
rect 27905 6069 27939 6103
rect 34161 6069 34195 6103
rect 39681 6069 39715 6103
rect 47869 6069 47903 6103
rect 52193 6069 52227 6103
rect 55781 6069 55815 6103
rect 56333 6069 56367 6103
rect 56885 6069 56919 6103
rect 2421 5865 2455 5899
rect 25881 5865 25915 5899
rect 27169 5865 27203 5899
rect 31401 5865 31435 5899
rect 34069 5865 34103 5899
rect 37565 5865 37599 5899
rect 42165 5865 42199 5899
rect 46765 5865 46799 5899
rect 50537 5865 50571 5899
rect 51549 5865 51583 5899
rect 56057 5865 56091 5899
rect 56609 5865 56643 5899
rect 57161 5865 57195 5899
rect 58357 5865 58391 5899
rect 31677 5797 31711 5831
rect 44281 5797 44315 5831
rect 45385 5797 45419 5831
rect 48329 5797 48363 5831
rect 50629 5797 50663 5831
rect 55505 5797 55539 5831
rect 26525 5729 26559 5763
rect 31769 5729 31803 5763
rect 32597 5729 32631 5763
rect 33149 5729 33183 5763
rect 36277 5729 36311 5763
rect 36369 5729 36403 5763
rect 37013 5729 37047 5763
rect 37105 5729 37139 5763
rect 41245 5729 41279 5763
rect 41613 5729 41647 5763
rect 41705 5729 41739 5763
rect 43361 5729 43395 5763
rect 45293 5729 45327 5763
rect 48697 5729 48731 5763
rect 52193 5729 52227 5763
rect 53113 5729 53147 5763
rect 54125 5729 54159 5763
rect 57713 5729 57747 5763
rect 1869 5661 1903 5695
rect 26065 5661 26099 5695
rect 26157 5661 26191 5695
rect 27350 5661 27384 5695
rect 27721 5661 27755 5695
rect 27813 5661 27847 5695
rect 28273 5661 28307 5695
rect 28457 5661 28491 5695
rect 28733 5661 28767 5695
rect 30021 5661 30055 5695
rect 30113 5661 30147 5695
rect 30205 5661 30239 5695
rect 30389 5661 30423 5695
rect 31585 5661 31619 5695
rect 31861 5661 31895 5695
rect 33333 5661 33367 5695
rect 33425 5661 33459 5695
rect 35265 5661 35299 5695
rect 35967 5661 36001 5695
rect 38025 5661 38059 5695
rect 38183 5661 38217 5695
rect 38301 5661 38335 5695
rect 38485 5661 38519 5695
rect 39313 5661 39347 5695
rect 41337 5661 41371 5695
rect 43269 5661 43303 5695
rect 44005 5661 44039 5695
rect 45201 5661 45235 5695
rect 46949 5661 46983 5695
rect 47041 5661 47075 5695
rect 47317 5661 47351 5695
rect 47409 5661 47443 5695
rect 48053 5661 48087 5695
rect 48605 5661 48639 5695
rect 49341 5661 49375 5695
rect 50997 5661 51031 5695
rect 52469 5661 52503 5695
rect 53389 5661 53423 5695
rect 54217 5661 54251 5695
rect 54861 5661 54895 5695
rect 25421 5593 25455 5627
rect 26433 5593 26467 5627
rect 37197 5593 37231 5627
rect 38393 5593 38427 5627
rect 39221 5593 39255 5627
rect 44281 5593 44315 5627
rect 45661 5593 45695 5627
rect 47133 5593 47167 5627
rect 1685 5525 1719 5559
rect 27353 5525 27387 5559
rect 28641 5525 28675 5559
rect 29745 5525 29779 5559
rect 35081 5525 35115 5559
rect 35817 5525 35851 5559
rect 38669 5525 38703 5559
rect 40141 5525 40175 5559
rect 41061 5525 41095 5559
rect 42901 5525 42935 5559
rect 44097 5525 44131 5559
rect 45569 5525 45603 5559
rect 46121 5525 46155 5559
rect 54861 5525 54895 5559
rect 26157 5321 26191 5355
rect 27353 5321 27387 5355
rect 28933 5321 28967 5355
rect 29101 5321 29135 5355
rect 30113 5321 30147 5355
rect 31769 5321 31803 5355
rect 32781 5321 32815 5355
rect 33793 5321 33827 5355
rect 36277 5321 36311 5355
rect 41429 5321 41463 5355
rect 45661 5321 45695 5355
rect 46857 5321 46891 5355
rect 48421 5321 48455 5355
rect 50261 5321 50295 5355
rect 51457 5321 51491 5355
rect 53205 5321 53239 5355
rect 55965 5321 55999 5355
rect 28733 5253 28767 5287
rect 36829 5253 36863 5287
rect 40325 5253 40359 5287
rect 42625 5253 42659 5287
rect 47869 5253 47903 5287
rect 53849 5253 53883 5287
rect 54953 5253 54987 5287
rect 55505 5253 55539 5287
rect 26433 5185 26467 5219
rect 27445 5185 27479 5219
rect 27629 5185 27663 5219
rect 27813 5185 27847 5219
rect 29561 5185 29595 5219
rect 29653 5185 29687 5219
rect 29837 5185 29871 5219
rect 29929 5185 29963 5219
rect 31125 5185 31159 5219
rect 31309 5185 31343 5219
rect 31401 5185 31435 5219
rect 31493 5185 31527 5219
rect 33701 5185 33735 5219
rect 33885 5185 33919 5219
rect 37749 5185 37783 5219
rect 37841 5185 37875 5219
rect 37933 5185 37967 5219
rect 38117 5185 38151 5219
rect 41521 5185 41555 5219
rect 44649 5185 44683 5219
rect 47041 5185 47075 5219
rect 48881 5185 48915 5219
rect 49341 5185 49375 5219
rect 51641 5185 51675 5219
rect 52377 5185 52411 5219
rect 53297 5185 53331 5219
rect 54585 5185 54619 5219
rect 57069 5185 57103 5219
rect 27353 5117 27387 5151
rect 33241 5117 33275 5151
rect 34529 5117 34563 5151
rect 34805 5117 34839 5151
rect 38577 5117 38611 5151
rect 40601 5117 40635 5151
rect 41705 5117 41739 5151
rect 44373 5117 44407 5151
rect 49525 5117 49559 5151
rect 27537 5049 27571 5083
rect 32873 5049 32907 5083
rect 52193 5049 52227 5083
rect 28917 4981 28951 5015
rect 30573 4981 30607 5015
rect 37565 4981 37599 5015
rect 41061 4981 41095 5015
rect 45109 4981 45143 5015
rect 46305 4981 46339 5015
rect 48789 4981 48823 5015
rect 50813 4981 50847 5015
rect 56517 4981 56551 5015
rect 26249 4777 26283 4811
rect 26709 4777 26743 4811
rect 27261 4777 27295 4811
rect 27813 4777 27847 4811
rect 29101 4777 29135 4811
rect 30113 4777 30147 4811
rect 31033 4777 31067 4811
rect 32505 4777 32539 4811
rect 33977 4777 34011 4811
rect 38301 4777 38335 4811
rect 39129 4777 39163 4811
rect 45845 4777 45879 4811
rect 47409 4777 47443 4811
rect 50353 4777 50387 4811
rect 51549 4777 51583 4811
rect 52745 4777 52779 4811
rect 54217 4777 54251 4811
rect 56057 4777 56091 4811
rect 56609 4777 56643 4811
rect 28089 4709 28123 4743
rect 29745 4709 29779 4743
rect 31861 4709 31895 4743
rect 34345 4709 34379 4743
rect 43729 4709 43763 4743
rect 49157 4709 49191 4743
rect 53573 4709 53607 4743
rect 55505 4709 55539 4743
rect 28181 4641 28215 4675
rect 30205 4641 30239 4675
rect 37841 4641 37875 4675
rect 45201 4641 45235 4675
rect 50905 4641 50939 4675
rect 54769 4641 54803 4675
rect 27997 4573 28031 4607
rect 28273 4573 28307 4607
rect 28457 4573 28491 4607
rect 29009 4573 29043 4607
rect 29193 4573 29227 4607
rect 29929 4573 29963 4607
rect 32413 4573 32447 4607
rect 32873 4573 32907 4607
rect 38301 4573 38335 4607
rect 39037 4573 39071 4607
rect 39221 4573 39255 4607
rect 41981 4573 42015 4607
rect 42901 4573 42935 4607
rect 46949 4573 46983 4607
rect 50721 4573 50755 4607
rect 53389 4573 53423 4607
rect 30941 4505 30975 4539
rect 34989 4505 35023 4539
rect 35357 4505 35391 4539
rect 35817 4505 35851 4539
rect 37565 4505 37599 4539
rect 42625 4505 42659 4539
rect 43453 4505 43487 4539
rect 44281 4505 44315 4539
rect 47961 4505 47995 4539
rect 50813 4505 50847 4539
rect 52469 4505 52503 4539
rect 33793 4437 33827 4471
rect 33977 4437 34011 4471
rect 40693 4437 40727 4471
rect 46305 4437 46339 4471
rect 48513 4437 48547 4471
rect 49617 4437 49651 4471
rect 33333 4233 33367 4267
rect 34069 4233 34103 4267
rect 34161 4233 34195 4267
rect 53849 4233 53883 4267
rect 54861 4233 54895 4267
rect 29101 4165 29135 4199
rect 31309 4165 31343 4199
rect 32413 4165 32447 4199
rect 34253 4165 34287 4199
rect 36645 4165 36679 4199
rect 41981 4165 42015 4199
rect 45010 4165 45044 4199
rect 48145 4165 48179 4199
rect 48973 4165 49007 4199
rect 52193 4165 52227 4199
rect 53113 4165 53147 4199
rect 53297 4165 53331 4199
rect 28181 4097 28215 4131
rect 28365 4097 28399 4131
rect 28457 4097 28491 4131
rect 30205 4097 30239 4131
rect 30665 4097 30699 4131
rect 31677 4097 31711 4131
rect 32321 4097 32355 4131
rect 32505 4097 32539 4131
rect 32689 4097 32723 4131
rect 33885 4097 33919 4131
rect 42625 4097 42659 4131
rect 43269 4097 43303 4131
rect 45293 4097 45327 4131
rect 45753 4097 45787 4131
rect 47225 4097 47259 4131
rect 48237 4097 48271 4131
rect 49525 4097 49559 4131
rect 50721 4097 50755 4131
rect 27997 4029 28031 4063
rect 34897 4029 34931 4063
rect 36921 4029 36955 4063
rect 37473 4029 37507 4063
rect 37749 4029 37783 4063
rect 39773 4029 39807 4063
rect 40049 4029 40083 4063
rect 48421 4029 48455 4063
rect 52929 4029 52963 4063
rect 55965 4029 55999 4063
rect 28273 3961 28307 3995
rect 29745 3961 29779 3995
rect 34437 3961 34471 3995
rect 41521 3961 41555 3995
rect 46305 3961 46339 3995
rect 47777 3961 47811 3995
rect 50169 3961 50203 3995
rect 30113 3893 30147 3927
rect 39221 3893 39255 3927
rect 47041 3893 47075 3927
rect 51181 3893 51215 3927
rect 54309 3893 54343 3927
rect 55413 3893 55447 3927
rect 28549 3689 28583 3723
rect 29745 3689 29779 3723
rect 30941 3689 30975 3723
rect 31309 3689 31343 3723
rect 31861 3689 31895 3723
rect 33609 3689 33643 3723
rect 33793 3689 33827 3723
rect 38669 3689 38703 3723
rect 47593 3689 47627 3723
rect 49341 3689 49375 3723
rect 53665 3689 53699 3723
rect 54677 3689 54711 3723
rect 55505 3689 55539 3723
rect 34989 3621 35023 3655
rect 40325 3621 40359 3655
rect 44281 3621 44315 3655
rect 48053 3621 48087 3655
rect 49249 3621 49283 3655
rect 54125 3621 54159 3655
rect 29929 3553 29963 3587
rect 30389 3553 30423 3587
rect 34253 3553 34287 3587
rect 37657 3553 37691 3587
rect 40969 3553 41003 3587
rect 41245 3553 41279 3587
rect 42993 3553 43027 3587
rect 45845 3553 45879 3587
rect 46121 3553 46155 3587
rect 30021 3485 30055 3519
rect 30849 3485 30883 3519
rect 32413 3485 32447 3519
rect 32609 3485 32643 3519
rect 33793 3485 33827 3519
rect 34161 3485 34195 3519
rect 35173 3485 35207 3519
rect 38485 3485 38519 3519
rect 40509 3485 40543 3519
rect 43545 3485 43579 3519
rect 48881 3485 48915 3519
rect 50353 3485 50387 3519
rect 52193 3485 52227 3519
rect 52653 3485 52687 3519
rect 32321 3417 32355 3451
rect 32781 3417 32815 3451
rect 35633 3417 35667 3451
rect 37381 3417 37415 3451
rect 39129 3417 39163 3451
rect 43729 3417 43763 3451
rect 45293 3349 45327 3383
rect 31033 3145 31067 3179
rect 37565 3145 37599 3179
rect 41337 3145 41371 3179
rect 41797 3145 41831 3179
rect 47777 3145 47811 3179
rect 48881 3145 48915 3179
rect 49525 3145 49559 3179
rect 52009 3145 52043 3179
rect 52929 3145 52963 3179
rect 53481 3145 53515 3179
rect 54125 3145 54159 3179
rect 54585 3145 54619 3179
rect 55229 3145 55263 3179
rect 58265 3145 58299 3179
rect 30205 3077 30239 3111
rect 30421 3077 30455 3111
rect 31493 3077 31527 3111
rect 32413 3077 32447 3111
rect 32827 3077 32861 3111
rect 35357 3077 35391 3111
rect 39037 3077 39071 3111
rect 42901 3077 42935 3111
rect 45385 3077 45419 3111
rect 48421 3077 48455 3111
rect 50169 3077 50203 3111
rect 50721 3077 50755 3111
rect 29193 3009 29227 3043
rect 33057 3009 33091 3043
rect 35633 3009 35667 3043
rect 36461 3009 36495 3043
rect 38761 3009 38795 3043
rect 41705 3009 41739 3043
rect 45109 3009 45143 3043
rect 51457 3009 51491 3043
rect 38025 2941 38059 2975
rect 40785 2941 40819 2975
rect 41889 2941 41923 2975
rect 42625 2941 42659 2975
rect 44649 2941 44683 2975
rect 47133 2941 47167 2975
rect 30573 2873 30607 2907
rect 31217 2873 31251 2907
rect 33885 2873 33919 2907
rect 36277 2873 36311 2907
rect 29745 2805 29779 2839
rect 30389 2805 30423 2839
rect 32781 2805 32815 2839
rect 12449 2601 12483 2635
rect 29193 2601 29227 2635
rect 30205 2601 30239 2635
rect 31125 2601 31159 2635
rect 36829 2601 36863 2635
rect 40877 2601 40911 2635
rect 43913 2601 43947 2635
rect 45293 2601 45327 2635
rect 46397 2601 46431 2635
rect 47041 2601 47075 2635
rect 48421 2601 48455 2635
rect 48881 2601 48915 2635
rect 51089 2601 51123 2635
rect 51641 2601 51675 2635
rect 52193 2601 52227 2635
rect 52929 2601 52963 2635
rect 53481 2601 53515 2635
rect 56977 2601 57011 2635
rect 2421 2533 2455 2567
rect 30757 2533 30791 2567
rect 32413 2533 32447 2567
rect 34069 2533 34103 2567
rect 35173 2533 35207 2567
rect 41889 2533 41923 2567
rect 45845 2533 45879 2567
rect 49433 2533 49467 2567
rect 5733 2465 5767 2499
rect 37473 2465 37507 2499
rect 41429 2465 41463 2499
rect 1869 2397 1903 2431
rect 6009 2397 6043 2431
rect 6561 2397 6595 2431
rect 11989 2397 12023 2431
rect 17141 2397 17175 2431
rect 22293 2397 22327 2431
rect 28089 2397 28123 2431
rect 30021 2397 30055 2431
rect 31217 2397 31251 2431
rect 32597 2397 32631 2431
rect 33333 2397 33367 2431
rect 33609 2397 33643 2431
rect 34161 2397 34195 2431
rect 35449 2397 35483 2431
rect 36277 2397 36311 2431
rect 40049 2397 40083 2431
rect 42073 2397 42107 2431
rect 50629 2397 50663 2431
rect 54033 2397 54067 2431
rect 56425 2397 56459 2431
rect 58081 2397 58115 2431
rect 39221 2329 39255 2363
rect 42625 2329 42659 2363
rect 47777 2329 47811 2363
rect 1685 2261 1719 2295
rect 11805 2261 11839 2295
rect 16957 2261 16991 2295
rect 17693 2261 17727 2295
rect 22109 2261 22143 2295
rect 22845 2261 22879 2295
rect 27905 2261 27939 2295
rect 28641 2261 28675 2295
rect 31769 2261 31803 2295
rect 36093 2261 36127 2295
rect 40233 2261 40267 2295
rect 50445 2261 50479 2295
rect 56241 2261 56275 2295
rect 58265 2261 58299 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 1673 57579 1731 57585
rect 1673 57545 1685 57579
rect 1719 57576 1731 57579
rect 2774 57576 2780 57588
rect 1719 57548 2780 57576
rect 1719 57545 1731 57548
rect 1673 57539 1731 57545
rect 2774 57536 2780 57548
rect 2832 57536 2838 57588
rect 3878 57536 3884 57588
rect 3936 57576 3942 57588
rect 4065 57579 4123 57585
rect 4065 57576 4077 57579
rect 3936 57548 4077 57576
rect 3936 57536 3942 57548
rect 4065 57545 4077 57548
rect 4111 57545 4123 57579
rect 4065 57539 4123 57545
rect 9674 57536 9680 57588
rect 9732 57576 9738 57588
rect 9861 57579 9919 57585
rect 9861 57576 9873 57579
rect 9732 57548 9873 57576
rect 9732 57536 9738 57548
rect 9861 57545 9873 57548
rect 9907 57545 9919 57579
rect 9861 57539 9919 57545
rect 15470 57536 15476 57588
rect 15528 57576 15534 57588
rect 15657 57579 15715 57585
rect 15657 57576 15669 57579
rect 15528 57548 15669 57576
rect 15528 57536 15534 57548
rect 15657 57545 15669 57548
rect 15703 57545 15715 57579
rect 15657 57539 15715 57545
rect 21266 57536 21272 57588
rect 21324 57576 21330 57588
rect 22097 57579 22155 57585
rect 22097 57576 22109 57579
rect 21324 57548 22109 57576
rect 21324 57536 21330 57548
rect 22097 57545 22109 57548
rect 22143 57545 22155 57579
rect 22097 57539 22155 57545
rect 26418 57536 26424 57588
rect 26476 57576 26482 57588
rect 27249 57579 27307 57585
rect 27249 57576 27261 57579
rect 26476 57548 27261 57576
rect 26476 57536 26482 57548
rect 27249 57545 27261 57548
rect 27295 57545 27307 57579
rect 27249 57539 27307 57545
rect 38010 57536 38016 57588
rect 38068 57576 38074 57588
rect 38289 57579 38347 57585
rect 38289 57576 38301 57579
rect 38068 57548 38301 57576
rect 38068 57536 38074 57548
rect 38289 57545 38301 57548
rect 38335 57545 38347 57579
rect 38289 57539 38347 57545
rect 43162 57536 43168 57588
rect 43220 57576 43226 57588
rect 43349 57579 43407 57585
rect 43349 57576 43361 57579
rect 43220 57548 43361 57576
rect 43220 57536 43226 57548
rect 43349 57545 43361 57548
rect 43395 57545 43407 57579
rect 43349 57539 43407 57545
rect 48958 57536 48964 57588
rect 49016 57576 49022 57588
rect 49145 57579 49203 57585
rect 49145 57576 49157 57579
rect 49016 57548 49157 57576
rect 49016 57536 49022 57548
rect 49145 57545 49157 57548
rect 49191 57545 49203 57579
rect 49145 57539 49203 57545
rect 54754 57536 54760 57588
rect 54812 57576 54818 57588
rect 55677 57579 55735 57585
rect 55677 57576 55689 57579
rect 54812 57548 55689 57576
rect 54812 57536 54818 57548
rect 55677 57545 55689 57548
rect 55723 57545 55735 57579
rect 58250 57576 58256 57588
rect 58211 57548 58256 57576
rect 55677 57539 55735 57545
rect 58250 57536 58256 57548
rect 58308 57536 58314 57588
rect 28718 57468 28724 57520
rect 28776 57508 28782 57520
rect 37553 57511 37611 57517
rect 37553 57508 37565 57511
rect 28776 57480 37565 57508
rect 28776 57468 28782 57480
rect 37553 57477 37565 57480
rect 37599 57508 37611 57511
rect 37599 57480 38148 57508
rect 37599 57477 37611 57480
rect 37553 57471 37611 57477
rect 1857 57443 1915 57449
rect 1857 57409 1869 57443
rect 1903 57440 1915 57443
rect 2314 57440 2320 57452
rect 1903 57412 2320 57440
rect 1903 57409 1915 57412
rect 1857 57403 1915 57409
rect 2314 57400 2320 57412
rect 2372 57400 2378 57452
rect 4249 57443 4307 57449
rect 4249 57409 4261 57443
rect 4295 57440 4307 57443
rect 4706 57440 4712 57452
rect 4295 57412 4712 57440
rect 4295 57409 4307 57412
rect 4249 57403 4307 57409
rect 4706 57400 4712 57412
rect 4764 57400 4770 57452
rect 10042 57440 10048 57452
rect 10003 57412 10048 57440
rect 10042 57400 10048 57412
rect 10100 57440 10106 57452
rect 10505 57443 10563 57449
rect 10505 57440 10517 57443
rect 10100 57412 10517 57440
rect 10100 57400 10106 57412
rect 10505 57409 10517 57412
rect 10551 57409 10563 57443
rect 10505 57403 10563 57409
rect 15841 57443 15899 57449
rect 15841 57409 15853 57443
rect 15887 57440 15899 57443
rect 15930 57440 15936 57452
rect 15887 57412 15936 57440
rect 15887 57409 15899 57412
rect 15841 57403 15899 57409
rect 15930 57400 15936 57412
rect 15988 57400 15994 57452
rect 22281 57443 22339 57449
rect 22281 57409 22293 57443
rect 22327 57440 22339 57443
rect 22646 57440 22652 57452
rect 22327 57412 22652 57440
rect 22327 57409 22339 57412
rect 22281 57403 22339 57409
rect 22646 57400 22652 57412
rect 22704 57400 22710 57452
rect 27433 57443 27491 57449
rect 27433 57409 27445 57443
rect 27479 57440 27491 57443
rect 27982 57440 27988 57452
rect 27479 57412 27988 57440
rect 27479 57409 27491 57412
rect 27433 57403 27491 57409
rect 27982 57400 27988 57412
rect 28040 57400 28046 57452
rect 31757 57443 31815 57449
rect 31757 57409 31769 57443
rect 31803 57440 31815 57443
rect 32214 57440 32220 57452
rect 31803 57412 32220 57440
rect 31803 57409 31815 57412
rect 31757 57403 31815 57409
rect 32214 57400 32220 57412
rect 32272 57440 32278 57452
rect 38120 57449 38148 57480
rect 32309 57443 32367 57449
rect 32309 57440 32321 57443
rect 32272 57412 32321 57440
rect 32272 57400 32278 57412
rect 32309 57409 32321 57412
rect 32355 57409 32367 57443
rect 32309 57403 32367 57409
rect 38105 57443 38163 57449
rect 38105 57409 38117 57443
rect 38151 57409 38163 57443
rect 38105 57403 38163 57409
rect 43533 57443 43591 57449
rect 43533 57409 43545 57443
rect 43579 57440 43591 57443
rect 43714 57440 43720 57452
rect 43579 57412 43720 57440
rect 43579 57409 43591 57412
rect 43533 57403 43591 57409
rect 43714 57400 43720 57412
rect 43772 57400 43778 57452
rect 49234 57400 49240 57452
rect 49292 57440 49298 57452
rect 49329 57443 49387 57449
rect 49329 57440 49341 57443
rect 49292 57412 49341 57440
rect 49292 57400 49298 57412
rect 49329 57409 49341 57412
rect 49375 57409 49387 57443
rect 55490 57440 55496 57452
rect 55451 57412 55496 57440
rect 49329 57403 49387 57409
rect 55490 57400 55496 57412
rect 55548 57400 55554 57452
rect 57698 57400 57704 57452
rect 57756 57440 57762 57452
rect 58069 57443 58127 57449
rect 58069 57440 58081 57443
rect 57756 57412 58081 57440
rect 57756 57400 57762 57412
rect 58069 57409 58081 57412
rect 58115 57409 58127 57443
rect 58069 57403 58127 57409
rect 32030 57332 32036 57384
rect 32088 57372 32094 57384
rect 32493 57375 32551 57381
rect 32493 57372 32505 57375
rect 32088 57344 32505 57372
rect 32088 57332 32094 57344
rect 32493 57341 32505 57344
rect 32539 57341 32551 57375
rect 32493 57335 32551 57341
rect 2314 57236 2320 57248
rect 2275 57208 2320 57236
rect 2314 57196 2320 57208
rect 2372 57196 2378 57248
rect 4706 57236 4712 57248
rect 4667 57208 4712 57236
rect 4706 57196 4712 57208
rect 4764 57196 4770 57248
rect 22646 57196 22652 57248
rect 22704 57236 22710 57248
rect 22741 57239 22799 57245
rect 22741 57236 22753 57239
rect 22704 57208 22753 57236
rect 22704 57196 22710 57208
rect 22741 57205 22753 57208
rect 22787 57205 22799 57239
rect 27982 57236 27988 57248
rect 27943 57208 27988 57236
rect 22741 57199 22799 57205
rect 27982 57196 27988 57208
rect 28040 57196 28046 57248
rect 43714 57196 43720 57248
rect 43772 57236 43778 57248
rect 43993 57239 44051 57245
rect 43993 57236 44005 57239
rect 43772 57208 44005 57236
rect 43772 57196 43778 57208
rect 43993 57205 44005 57208
rect 44039 57205 44051 57239
rect 43993 57199 44051 57205
rect 57517 57239 57575 57245
rect 57517 57205 57529 57239
rect 57563 57236 57575 57239
rect 57698 57236 57704 57248
rect 57563 57208 57704 57236
rect 57563 57205 57575 57208
rect 57517 57199 57575 57205
rect 57698 57196 57704 57208
rect 57756 57196 57762 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 40402 56788 40408 56840
rect 40460 56828 40466 56840
rect 41141 56831 41199 56837
rect 41141 56828 41153 56831
rect 40460 56800 41153 56828
rect 40460 56788 40466 56800
rect 41141 56797 41153 56800
rect 41187 56828 41199 56831
rect 41785 56831 41843 56837
rect 41785 56828 41797 56831
rect 41187 56800 41797 56828
rect 41187 56797 41199 56800
rect 41141 56791 41199 56797
rect 41785 56797 41797 56800
rect 41831 56797 41843 56831
rect 41785 56791 41843 56797
rect 55490 56760 55496 56772
rect 41340 56732 55496 56760
rect 15930 56692 15936 56704
rect 15891 56664 15936 56692
rect 15930 56652 15936 56664
rect 15988 56652 15994 56704
rect 41340 56701 41368 56732
rect 55490 56720 55496 56732
rect 55548 56720 55554 56772
rect 41325 56695 41383 56701
rect 41325 56661 41337 56695
rect 41371 56661 41383 56695
rect 41325 56655 41383 56661
rect 49234 56652 49240 56704
rect 49292 56692 49298 56704
rect 49421 56695 49479 56701
rect 49421 56692 49433 56695
rect 49292 56664 49433 56692
rect 49292 56652 49298 56664
rect 49421 56661 49433 56664
rect 49467 56661 49479 56695
rect 49421 56655 49479 56661
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 58069 54655 58127 54661
rect 58069 54652 58081 54655
rect 57532 54624 58081 54652
rect 57330 54476 57336 54528
rect 57388 54516 57394 54528
rect 57532 54525 57560 54624
rect 58069 54621 58081 54624
rect 58115 54621 58127 54655
rect 58069 54615 58127 54621
rect 57517 54519 57575 54525
rect 57517 54516 57529 54519
rect 57388 54488 57529 54516
rect 57388 54476 57394 54488
rect 57517 54485 57529 54488
rect 57563 54485 57575 54519
rect 58250 54516 58256 54528
rect 58211 54488 58256 54516
rect 57517 54479 57575 54485
rect 58250 54476 58256 54488
rect 58308 54476 58314 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1857 53567 1915 53573
rect 1857 53533 1869 53567
rect 1903 53564 1915 53567
rect 1903 53536 2452 53564
rect 1903 53533 1915 53536
rect 1857 53527 1915 53533
rect 2424 53440 2452 53536
rect 1670 53428 1676 53440
rect 1631 53400 1676 53428
rect 1670 53388 1676 53400
rect 1728 53388 1734 53440
rect 2406 53428 2412 53440
rect 2367 53400 2412 53428
rect 2406 53388 2412 53400
rect 2464 53388 2470 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 57790 48696 57796 48748
rect 57848 48736 57854 48748
rect 58069 48739 58127 48745
rect 58069 48736 58081 48739
rect 57848 48708 58081 48736
rect 57848 48696 57854 48708
rect 58069 48705 58081 48708
rect 58115 48705 58127 48739
rect 58069 48699 58127 48705
rect 57517 48535 57575 48541
rect 57517 48501 57529 48535
rect 57563 48532 57575 48535
rect 57790 48532 57796 48544
rect 57563 48504 57796 48532
rect 57563 48501 57575 48504
rect 57517 48495 57575 48501
rect 57790 48492 57796 48504
rect 57848 48492 57854 48544
rect 58250 48532 58256 48544
rect 58211 48504 58256 48532
rect 58250 48492 58256 48504
rect 58308 48492 58314 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1670 47172 1676 47184
rect 1631 47144 1676 47172
rect 1670 47132 1676 47144
rect 1728 47132 1734 47184
rect 1857 47039 1915 47045
rect 1857 47005 1869 47039
rect 1903 47005 1915 47039
rect 1857 46999 1915 47005
rect 1872 46968 1900 46999
rect 2409 46971 2467 46977
rect 2409 46968 2421 46971
rect 1872 46940 2421 46968
rect 2409 46937 2421 46940
rect 2455 46968 2467 46971
rect 2498 46968 2504 46980
rect 2455 46940 2504 46968
rect 2455 46937 2467 46940
rect 2409 46931 2467 46937
rect 2498 46928 2504 46940
rect 2556 46928 2562 46980
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 58069 42687 58127 42693
rect 58069 42684 58081 42687
rect 57532 42656 58081 42684
rect 57532 42560 57560 42656
rect 58069 42653 58081 42656
rect 58115 42653 58127 42687
rect 58069 42647 58127 42653
rect 57514 42548 57520 42560
rect 57475 42520 57520 42548
rect 57514 42508 57520 42520
rect 57572 42508 57578 42560
rect 58250 42548 58256 42560
rect 58211 42520 58256 42548
rect 58250 42508 58256 42520
rect 58308 42508 58314 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1854 41120 1860 41132
rect 1815 41092 1860 41120
rect 1854 41080 1860 41092
rect 1912 41120 1918 41132
rect 2317 41123 2375 41129
rect 2317 41120 2329 41123
rect 1912 41092 2329 41120
rect 1912 41080 1918 41092
rect 2317 41089 2329 41092
rect 2363 41089 2375 41123
rect 2317 41083 2375 41089
rect 1670 40916 1676 40928
rect 1631 40888 1676 40916
rect 1670 40876 1676 40888
rect 1728 40876 1734 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 57974 37204 57980 37256
rect 58032 37244 58038 37256
rect 58069 37247 58127 37253
rect 58069 37244 58081 37247
rect 58032 37216 58081 37244
rect 58032 37204 58038 37216
rect 58069 37213 58081 37216
rect 58115 37213 58127 37247
rect 58069 37207 58127 37213
rect 58250 37108 58256 37120
rect 58211 37080 58256 37108
rect 58250 37068 58256 37080
rect 58308 37068 58314 37120
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1857 35683 1915 35689
rect 1857 35649 1869 35683
rect 1903 35680 1915 35683
rect 1946 35680 1952 35692
rect 1903 35652 1952 35680
rect 1903 35649 1915 35652
rect 1857 35643 1915 35649
rect 1946 35640 1952 35652
rect 2004 35680 2010 35692
rect 2317 35683 2375 35689
rect 2317 35680 2329 35683
rect 2004 35652 2329 35680
rect 2004 35640 2010 35652
rect 2317 35649 2329 35652
rect 2363 35649 2375 35683
rect 2317 35643 2375 35649
rect 1670 35476 1676 35488
rect 1631 35448 1676 35476
rect 1670 35436 1676 35448
rect 1728 35436 1734 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 44818 31328 44824 31340
rect 44779 31300 44824 31328
rect 44818 31288 44824 31300
rect 44876 31288 44882 31340
rect 44910 31288 44916 31340
rect 44968 31328 44974 31340
rect 45189 31331 45247 31337
rect 45189 31328 45201 31331
rect 44968 31300 45201 31328
rect 44968 31288 44974 31300
rect 45189 31297 45201 31300
rect 45235 31297 45247 31331
rect 46750 31328 46756 31340
rect 46711 31300 46756 31328
rect 45189 31291 45247 31297
rect 46750 31288 46756 31300
rect 46808 31288 46814 31340
rect 47026 31328 47032 31340
rect 46987 31300 47032 31328
rect 47026 31288 47032 31300
rect 47084 31288 47090 31340
rect 4706 31084 4712 31136
rect 4764 31124 4770 31136
rect 44269 31127 44327 31133
rect 44269 31124 44281 31127
rect 4764 31096 44281 31124
rect 4764 31084 4770 31096
rect 44269 31093 44281 31096
rect 44315 31093 44327 31127
rect 46934 31124 46940 31136
rect 46895 31096 46940 31124
rect 44269 31087 44327 31093
rect 46934 31084 46940 31096
rect 46992 31084 46998 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 48406 30744 48412 30796
rect 48464 30784 48470 30796
rect 49234 30784 49240 30796
rect 48464 30756 48509 30784
rect 49195 30756 49240 30784
rect 48464 30744 48470 30756
rect 49234 30744 49240 30756
rect 49292 30744 49298 30796
rect 48320 30728 48372 30734
rect 46290 30716 46296 30728
rect 46251 30688 46296 30716
rect 46290 30676 46296 30688
rect 46348 30676 46354 30728
rect 46934 30716 46940 30728
rect 46895 30688 46940 30716
rect 46934 30676 46940 30688
rect 46992 30676 46998 30728
rect 58069 30719 58127 30725
rect 58069 30685 58081 30719
rect 58115 30716 58127 30719
rect 58158 30716 58164 30728
rect 58115 30688 58164 30716
rect 58115 30685 58127 30688
rect 58069 30679 58127 30685
rect 58158 30676 58164 30688
rect 58216 30676 58222 30728
rect 48320 30670 48372 30676
rect 2406 30608 2412 30660
rect 2464 30648 2470 30660
rect 45741 30651 45799 30657
rect 45741 30648 45753 30651
rect 2464 30620 45753 30648
rect 2464 30608 2470 30620
rect 45741 30617 45753 30620
rect 45787 30617 45799 30651
rect 45741 30611 45799 30617
rect 58250 30580 58256 30592
rect 58211 30552 58256 30580
rect 58250 30540 58256 30552
rect 58308 30540 58314 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 46201 30379 46259 30385
rect 46201 30345 46213 30379
rect 46247 30376 46259 30379
rect 46750 30376 46756 30388
rect 46247 30348 46756 30376
rect 46247 30345 46259 30348
rect 46201 30339 46259 30345
rect 46750 30336 46756 30348
rect 46808 30336 46814 30388
rect 44818 30308 44824 30320
rect 44779 30280 44824 30308
rect 44818 30268 44824 30280
rect 44876 30268 44882 30320
rect 46109 30311 46167 30317
rect 46109 30277 46121 30311
rect 46155 30308 46167 30311
rect 46290 30308 46296 30320
rect 46155 30280 46296 30308
rect 46155 30277 46167 30280
rect 46109 30271 46167 30277
rect 45281 30175 45339 30181
rect 45281 30141 45293 30175
rect 45327 30172 45339 30175
rect 46124 30172 46152 30271
rect 46290 30268 46296 30280
rect 46348 30268 46354 30320
rect 46569 30311 46627 30317
rect 46569 30277 46581 30311
rect 46615 30308 46627 30311
rect 48314 30308 48320 30320
rect 46615 30280 48320 30308
rect 46615 30277 46627 30280
rect 46569 30271 46627 30277
rect 48314 30268 48320 30280
rect 48372 30308 48378 30320
rect 49510 30308 49516 30320
rect 48372 30280 49516 30308
rect 48372 30268 48378 30280
rect 49510 30268 49516 30280
rect 49568 30308 49574 30320
rect 49789 30311 49847 30317
rect 49789 30308 49801 30311
rect 49568 30280 49801 30308
rect 49568 30268 49574 30280
rect 49789 30277 49801 30280
rect 49835 30277 49847 30311
rect 49789 30271 49847 30277
rect 46382 30240 46388 30252
rect 46343 30212 46388 30240
rect 46382 30200 46388 30212
rect 46440 30200 46446 30252
rect 49234 30200 49240 30252
rect 49292 30240 49298 30252
rect 49605 30243 49663 30249
rect 49605 30240 49617 30243
rect 49292 30212 49617 30240
rect 49292 30200 49298 30212
rect 49605 30209 49617 30212
rect 49651 30209 49663 30243
rect 49605 30203 49663 30209
rect 45327 30144 46152 30172
rect 45327 30141 45339 30144
rect 45281 30135 45339 30141
rect 44910 30064 44916 30116
rect 44968 30104 44974 30116
rect 45097 30107 45155 30113
rect 45097 30104 45109 30107
rect 44968 30076 45109 30104
rect 44968 30064 44974 30076
rect 45097 30073 45109 30076
rect 45143 30073 45155 30107
rect 45097 30067 45155 30073
rect 49418 30036 49424 30048
rect 49379 30008 49424 30036
rect 49418 29996 49424 30008
rect 49476 29996 49482 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 46750 29832 46756 29844
rect 46711 29804 46756 29832
rect 46750 29792 46756 29804
rect 46808 29792 46814 29844
rect 47026 29792 47032 29844
rect 47084 29832 47090 29844
rect 47305 29835 47363 29841
rect 47305 29832 47317 29835
rect 47084 29804 47317 29832
rect 47084 29792 47090 29804
rect 47305 29801 47317 29804
rect 47351 29801 47363 29835
rect 47305 29795 47363 29801
rect 48406 29792 48412 29844
rect 48464 29832 48470 29844
rect 48777 29835 48835 29841
rect 48777 29832 48789 29835
rect 48464 29804 48789 29832
rect 48464 29792 48470 29804
rect 48777 29801 48789 29804
rect 48823 29801 48835 29835
rect 48777 29795 48835 29801
rect 46382 29724 46388 29776
rect 46440 29764 46446 29776
rect 48130 29764 48136 29776
rect 46440 29736 47256 29764
rect 48091 29736 48136 29764
rect 46440 29724 46446 29736
rect 44726 29656 44732 29708
rect 44784 29696 44790 29708
rect 45649 29699 45707 29705
rect 45649 29696 45661 29699
rect 44784 29668 45661 29696
rect 44784 29656 44790 29668
rect 45649 29665 45661 29668
rect 45695 29665 45707 29699
rect 45649 29659 45707 29665
rect 45833 29699 45891 29705
rect 45833 29665 45845 29699
rect 45879 29696 45891 29699
rect 46106 29696 46112 29708
rect 45879 29668 46112 29696
rect 45879 29665 45891 29668
rect 45833 29659 45891 29665
rect 46106 29656 46112 29668
rect 46164 29696 46170 29708
rect 46164 29668 46612 29696
rect 46164 29656 46170 29668
rect 1857 29631 1915 29637
rect 1857 29597 1869 29631
rect 1903 29628 1915 29631
rect 1903 29600 2452 29628
rect 1903 29597 1915 29600
rect 1857 29591 1915 29597
rect 2424 29504 2452 29600
rect 45462 29588 45468 29640
rect 45520 29628 45526 29640
rect 45557 29631 45615 29637
rect 45557 29628 45569 29631
rect 45520 29600 45569 29628
rect 45520 29588 45526 29600
rect 45557 29597 45569 29600
rect 45603 29597 45615 29631
rect 45557 29591 45615 29597
rect 46198 29588 46204 29640
rect 46256 29628 46262 29640
rect 46584 29637 46612 29668
rect 47228 29637 47256 29736
rect 48130 29724 48136 29736
rect 48188 29724 48194 29776
rect 48958 29764 48964 29776
rect 48919 29736 48964 29764
rect 48958 29724 48964 29736
rect 49016 29724 49022 29776
rect 51997 29767 52055 29773
rect 51997 29733 52009 29767
rect 52043 29764 52055 29767
rect 57514 29764 57520 29776
rect 52043 29736 57520 29764
rect 52043 29733 52055 29736
rect 51997 29727 52055 29733
rect 57514 29724 57520 29736
rect 57572 29724 57578 29776
rect 48317 29699 48375 29705
rect 48317 29665 48329 29699
rect 48363 29696 48375 29699
rect 49234 29696 49240 29708
rect 48363 29668 49240 29696
rect 48363 29665 48375 29668
rect 48317 29659 48375 29665
rect 49234 29656 49240 29668
rect 49292 29656 49298 29708
rect 50893 29699 50951 29705
rect 50893 29665 50905 29699
rect 50939 29696 50951 29699
rect 51537 29699 51595 29705
rect 51537 29696 51549 29699
rect 50939 29668 51549 29696
rect 50939 29665 50951 29668
rect 50893 29659 50951 29665
rect 51537 29665 51549 29668
rect 51583 29665 51595 29699
rect 51537 29659 51595 29665
rect 46293 29631 46351 29637
rect 46293 29628 46305 29631
rect 46256 29600 46305 29628
rect 46256 29588 46262 29600
rect 46293 29597 46305 29600
rect 46339 29597 46351 29631
rect 46293 29591 46351 29597
rect 46569 29631 46627 29637
rect 46569 29597 46581 29631
rect 46615 29597 46627 29631
rect 46569 29591 46627 29597
rect 47213 29631 47271 29637
rect 47213 29597 47225 29631
rect 47259 29597 47271 29631
rect 47213 29591 47271 29597
rect 50801 29631 50859 29637
rect 50801 29597 50813 29631
rect 50847 29597 50859 29631
rect 50982 29628 50988 29640
rect 50943 29600 50988 29628
rect 50801 29591 50859 29597
rect 47857 29563 47915 29569
rect 47857 29529 47869 29563
rect 47903 29560 47915 29563
rect 47946 29560 47952 29572
rect 47903 29532 47952 29560
rect 47903 29529 47915 29532
rect 47857 29523 47915 29529
rect 47946 29520 47952 29532
rect 48004 29520 48010 29572
rect 50816 29560 50844 29591
rect 50982 29588 50988 29600
rect 51040 29588 51046 29640
rect 51629 29631 51687 29637
rect 51629 29597 51641 29631
rect 51675 29628 51687 29631
rect 51810 29628 51816 29640
rect 51675 29600 51816 29628
rect 51675 29597 51687 29600
rect 51629 29591 51687 29597
rect 51810 29588 51816 29600
rect 51868 29588 51874 29640
rect 50816 29532 51028 29560
rect 51000 29504 51028 29532
rect 1670 29492 1676 29504
rect 1631 29464 1676 29492
rect 1670 29452 1676 29464
rect 1728 29452 1734 29504
rect 2406 29492 2412 29504
rect 2367 29464 2412 29492
rect 2406 29452 2412 29464
rect 2464 29452 2470 29504
rect 45186 29492 45192 29504
rect 45147 29464 45192 29492
rect 45186 29452 45192 29464
rect 45244 29452 45250 29504
rect 46385 29495 46443 29501
rect 46385 29461 46397 29495
rect 46431 29492 46443 29495
rect 47210 29492 47216 29504
rect 46431 29464 47216 29492
rect 46431 29461 46443 29464
rect 46385 29455 46443 29461
rect 47210 29452 47216 29464
rect 47268 29452 47274 29504
rect 50982 29452 50988 29504
rect 51040 29452 51046 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 44818 29248 44824 29300
rect 44876 29288 44882 29300
rect 45281 29291 45339 29297
rect 45281 29288 45293 29291
rect 44876 29260 45293 29288
rect 44876 29248 44882 29260
rect 45281 29257 45293 29260
rect 45327 29257 45339 29291
rect 45281 29251 45339 29257
rect 46106 29248 46112 29300
rect 46164 29297 46170 29300
rect 46164 29291 46183 29297
rect 46171 29257 46183 29291
rect 46164 29251 46183 29257
rect 46293 29291 46351 29297
rect 46293 29257 46305 29291
rect 46339 29288 46351 29291
rect 46382 29288 46388 29300
rect 46339 29260 46388 29288
rect 46339 29257 46351 29260
rect 46293 29251 46351 29257
rect 46164 29248 46170 29251
rect 46382 29248 46388 29260
rect 46440 29248 46446 29300
rect 49602 29248 49608 29300
rect 49660 29288 49666 29300
rect 51810 29288 51816 29300
rect 49660 29260 50384 29288
rect 51771 29260 51816 29288
rect 49660 29248 49666 29260
rect 45925 29223 45983 29229
rect 45925 29189 45937 29223
rect 45971 29189 45983 29223
rect 45925 29183 45983 29189
rect 44637 29155 44695 29161
rect 44637 29121 44649 29155
rect 44683 29152 44695 29155
rect 44818 29152 44824 29164
rect 44683 29124 44824 29152
rect 44683 29121 44695 29124
rect 44637 29115 44695 29121
rect 44818 29112 44824 29124
rect 44876 29152 44882 29164
rect 45462 29152 45468 29164
rect 44876 29124 45468 29152
rect 44876 29112 44882 29124
rect 45462 29112 45468 29124
rect 45520 29112 45526 29164
rect 45940 29152 45968 29183
rect 46753 29155 46811 29161
rect 46753 29152 46765 29155
rect 45940 29124 46765 29152
rect 46753 29121 46765 29124
rect 46799 29152 46811 29155
rect 47210 29152 47216 29164
rect 46799 29124 47216 29152
rect 46799 29121 46811 29124
rect 46753 29115 46811 29121
rect 47210 29112 47216 29124
rect 47268 29112 47274 29164
rect 47946 29152 47952 29164
rect 47907 29124 47952 29152
rect 47946 29112 47952 29124
rect 48004 29112 48010 29164
rect 49234 29152 49240 29164
rect 49195 29124 49240 29152
rect 49234 29112 49240 29124
rect 49292 29112 49298 29164
rect 49510 29112 49516 29164
rect 49568 29152 49574 29164
rect 49697 29155 49755 29161
rect 49697 29152 49709 29155
rect 49568 29124 49709 29152
rect 49568 29112 49574 29124
rect 49697 29121 49709 29124
rect 49743 29121 49755 29155
rect 49697 29115 49755 29121
rect 49786 29112 49792 29164
rect 49844 29152 49850 29164
rect 50356 29161 50384 29260
rect 51810 29248 51816 29260
rect 51868 29248 51874 29300
rect 50890 29180 50896 29232
rect 50948 29220 50954 29232
rect 51629 29223 51687 29229
rect 51629 29220 51641 29223
rect 50948 29192 51641 29220
rect 50948 29180 50954 29192
rect 51629 29189 51641 29192
rect 51675 29189 51687 29223
rect 51629 29183 51687 29189
rect 49973 29155 50031 29161
rect 49973 29152 49985 29155
rect 49844 29124 49985 29152
rect 49844 29112 49850 29124
rect 49973 29121 49985 29124
rect 50019 29121 50031 29155
rect 49973 29115 50031 29121
rect 50341 29155 50399 29161
rect 50341 29121 50353 29155
rect 50387 29121 50399 29155
rect 50341 29115 50399 29121
rect 50709 29155 50767 29161
rect 50709 29121 50721 29155
rect 50755 29121 50767 29155
rect 50709 29115 50767 29121
rect 44726 29084 44732 29096
rect 44687 29056 44732 29084
rect 44726 29044 44732 29056
rect 44784 29044 44790 29096
rect 48409 29087 48467 29093
rect 48409 29053 48421 29087
rect 48455 29084 48467 29087
rect 48958 29084 48964 29096
rect 48455 29056 48964 29084
rect 48455 29053 48467 29056
rect 48409 29047 48467 29053
rect 48958 29044 48964 29056
rect 49016 29084 49022 29096
rect 49326 29084 49332 29096
rect 49016 29056 49332 29084
rect 49016 29044 49022 29056
rect 49326 29044 49332 29056
rect 49384 29084 49390 29096
rect 50724 29084 50752 29115
rect 51166 29112 51172 29164
rect 51224 29152 51230 29164
rect 51445 29155 51503 29161
rect 51445 29152 51457 29155
rect 51224 29124 51457 29152
rect 51224 29112 51230 29124
rect 51445 29121 51457 29124
rect 51491 29121 51503 29155
rect 51445 29115 51503 29121
rect 53837 29155 53895 29161
rect 53837 29121 53849 29155
rect 53883 29152 53895 29155
rect 54110 29152 54116 29164
rect 53883 29124 54116 29152
rect 53883 29121 53895 29124
rect 53837 29115 53895 29121
rect 54110 29112 54116 29124
rect 54168 29112 54174 29164
rect 54481 29155 54539 29161
rect 54481 29121 54493 29155
rect 54527 29152 54539 29155
rect 55214 29152 55220 29164
rect 54527 29124 55220 29152
rect 54527 29121 54539 29124
rect 54481 29115 54539 29121
rect 55214 29112 55220 29124
rect 55272 29112 55278 29164
rect 49384 29056 50752 29084
rect 49384 29044 49390 29056
rect 1854 28976 1860 29028
rect 1912 29016 1918 29028
rect 53009 29019 53067 29025
rect 53009 29016 53021 29019
rect 1912 28988 53021 29016
rect 1912 28976 1918 28988
rect 53009 28985 53021 28988
rect 53055 28985 53067 29019
rect 53009 28979 53067 28985
rect 46109 28951 46167 28957
rect 46109 28917 46121 28951
rect 46155 28948 46167 28951
rect 46198 28948 46204 28960
rect 46155 28920 46204 28948
rect 46155 28917 46167 28920
rect 46109 28911 46167 28917
rect 46198 28908 46204 28920
rect 46256 28908 46262 28960
rect 46842 28948 46848 28960
rect 46803 28920 46848 28948
rect 46842 28908 46848 28920
rect 46900 28908 46906 28960
rect 47213 28951 47271 28957
rect 47213 28917 47225 28951
rect 47259 28948 47271 28951
rect 48130 28948 48136 28960
rect 47259 28920 48136 28948
rect 47259 28917 47271 28920
rect 47213 28911 47271 28917
rect 48130 28908 48136 28920
rect 48188 28908 48194 28960
rect 50982 28948 50988 28960
rect 50943 28920 50988 28948
rect 50982 28908 50988 28920
rect 51040 28908 51046 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 46198 28744 46204 28756
rect 46159 28716 46204 28744
rect 46198 28704 46204 28716
rect 46256 28704 46262 28756
rect 46753 28747 46811 28753
rect 46753 28713 46765 28747
rect 46799 28713 46811 28747
rect 47210 28744 47216 28756
rect 47171 28716 47216 28744
rect 46753 28707 46811 28713
rect 46014 28685 46020 28688
rect 45971 28679 46020 28685
rect 45971 28676 45983 28679
rect 45927 28648 45983 28676
rect 45971 28645 45983 28648
rect 46017 28645 46020 28679
rect 45971 28639 46020 28645
rect 46014 28636 46020 28639
rect 46072 28676 46078 28688
rect 46768 28676 46796 28707
rect 47210 28704 47216 28716
rect 47268 28704 47274 28756
rect 46072 28648 46796 28676
rect 49789 28679 49847 28685
rect 46072 28636 46078 28648
rect 49789 28645 49801 28679
rect 49835 28645 49847 28679
rect 49789 28639 49847 28645
rect 46109 28611 46167 28617
rect 46109 28577 46121 28611
rect 46155 28608 46167 28611
rect 46842 28608 46848 28620
rect 46155 28580 46848 28608
rect 46155 28577 46167 28580
rect 46109 28571 46167 28577
rect 46842 28568 46848 28580
rect 46900 28568 46906 28620
rect 49326 28608 49332 28620
rect 49252 28580 49332 28608
rect 45646 28500 45652 28552
rect 45704 28540 45710 28552
rect 49252 28549 49280 28580
rect 49326 28568 49332 28580
rect 49384 28568 49390 28620
rect 45833 28543 45891 28549
rect 45833 28540 45845 28543
rect 45704 28512 45845 28540
rect 45704 28500 45710 28512
rect 45833 28509 45845 28512
rect 45879 28509 45891 28543
rect 46293 28543 46351 28549
rect 46293 28542 46305 28543
rect 45833 28503 45891 28509
rect 46216 28514 46305 28542
rect 45002 28432 45008 28484
rect 45060 28472 45066 28484
rect 46216 28472 46244 28514
rect 46293 28509 46305 28514
rect 46339 28509 46351 28543
rect 46293 28503 46351 28509
rect 47029 28543 47087 28549
rect 47029 28509 47041 28543
rect 47075 28509 47087 28543
rect 47029 28503 47087 28509
rect 49237 28543 49295 28549
rect 49237 28509 49249 28543
rect 49283 28509 49295 28543
rect 49418 28540 49424 28552
rect 49379 28512 49424 28540
rect 49237 28503 49295 28509
rect 46753 28475 46811 28481
rect 46753 28472 46765 28475
rect 45060 28444 46765 28472
rect 45060 28432 45066 28444
rect 46753 28441 46765 28444
rect 46799 28441 46811 28475
rect 46753 28435 46811 28441
rect 45646 28364 45652 28416
rect 45704 28404 45710 28416
rect 46658 28404 46664 28416
rect 45704 28376 46664 28404
rect 45704 28364 45710 28376
rect 46658 28364 46664 28376
rect 46716 28404 46722 28416
rect 47044 28404 47072 28503
rect 49418 28500 49424 28512
rect 49476 28500 49482 28552
rect 49602 28540 49608 28552
rect 49563 28512 49608 28540
rect 49602 28500 49608 28512
rect 49660 28500 49666 28552
rect 49804 28540 49832 28639
rect 50798 28636 50804 28688
rect 50856 28676 50862 28688
rect 50856 28648 51672 28676
rect 50856 28636 50862 28648
rect 50709 28611 50767 28617
rect 50709 28577 50721 28611
rect 50755 28608 50767 28611
rect 50982 28608 50988 28620
rect 50755 28580 50988 28608
rect 50755 28577 50767 28580
rect 50709 28571 50767 28577
rect 50982 28568 50988 28580
rect 51040 28608 51046 28620
rect 51040 28580 51580 28608
rect 51040 28568 51046 28580
rect 50525 28543 50583 28549
rect 50525 28540 50537 28543
rect 49804 28512 50537 28540
rect 50525 28509 50537 28512
rect 50571 28509 50583 28543
rect 51350 28540 51356 28552
rect 51311 28512 51356 28540
rect 50525 28503 50583 28509
rect 51350 28500 51356 28512
rect 51408 28500 51414 28552
rect 51552 28549 51580 28580
rect 51537 28543 51595 28549
rect 51537 28509 51549 28543
rect 51583 28509 51595 28543
rect 51644 28540 51672 28648
rect 53926 28608 53932 28620
rect 53668 28580 53932 28608
rect 51905 28543 51963 28549
rect 51905 28540 51917 28543
rect 51644 28512 51917 28540
rect 51537 28503 51595 28509
rect 51905 28509 51917 28512
rect 51951 28509 51963 28543
rect 51905 28503 51963 28509
rect 52273 28543 52331 28549
rect 52273 28509 52285 28543
rect 52319 28509 52331 28543
rect 52914 28540 52920 28552
rect 52875 28512 52920 28540
rect 52273 28503 52331 28509
rect 49513 28475 49571 28481
rect 49513 28441 49525 28475
rect 49559 28472 49571 28475
rect 49786 28472 49792 28484
rect 49559 28444 49792 28472
rect 49559 28441 49571 28444
rect 49513 28435 49571 28441
rect 49786 28432 49792 28444
rect 49844 28432 49850 28484
rect 51166 28432 51172 28484
rect 51224 28472 51230 28484
rect 52288 28472 52316 28503
rect 52914 28500 52920 28512
rect 52972 28500 52978 28552
rect 53668 28549 53696 28580
rect 53926 28568 53932 28580
rect 53984 28568 53990 28620
rect 53653 28543 53711 28549
rect 53653 28509 53665 28543
rect 53699 28509 53711 28543
rect 53653 28503 53711 28509
rect 53742 28500 53748 28552
rect 53800 28540 53806 28552
rect 53837 28543 53895 28549
rect 53837 28540 53849 28543
rect 53800 28512 53849 28540
rect 53800 28500 53806 28512
rect 53837 28509 53849 28512
rect 53883 28509 53895 28543
rect 53837 28503 53895 28509
rect 56781 28543 56839 28549
rect 56781 28509 56793 28543
rect 56827 28509 56839 28543
rect 56781 28503 56839 28509
rect 56965 28543 57023 28549
rect 56965 28509 56977 28543
rect 57011 28540 57023 28543
rect 57146 28540 57152 28552
rect 57011 28512 57152 28540
rect 57011 28509 57023 28512
rect 56965 28503 57023 28509
rect 51224 28444 52316 28472
rect 56796 28472 56824 28503
rect 57146 28500 57152 28512
rect 57204 28500 57210 28552
rect 57238 28472 57244 28484
rect 56796 28444 57244 28472
rect 51224 28432 51230 28444
rect 57238 28432 57244 28444
rect 57296 28432 57302 28484
rect 46716 28376 47072 28404
rect 46716 28364 46722 28376
rect 50062 28364 50068 28416
rect 50120 28404 50126 28416
rect 50341 28407 50399 28413
rect 50341 28404 50353 28407
rect 50120 28376 50353 28404
rect 50120 28364 50126 28376
rect 50341 28373 50353 28376
rect 50387 28373 50399 28407
rect 53006 28404 53012 28416
rect 52967 28376 53012 28404
rect 50341 28367 50399 28373
rect 53006 28364 53012 28376
rect 53064 28364 53070 28416
rect 53834 28404 53840 28416
rect 53795 28376 53840 28404
rect 53834 28364 53840 28376
rect 53892 28364 53898 28416
rect 56962 28404 56968 28416
rect 56923 28376 56968 28404
rect 56962 28364 56968 28376
rect 57020 28364 57026 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 46569 28203 46627 28209
rect 46569 28169 46581 28203
rect 46615 28200 46627 28203
rect 46842 28200 46848 28212
rect 46615 28172 46848 28200
rect 46615 28169 46627 28172
rect 46569 28163 46627 28169
rect 46842 28160 46848 28172
rect 46900 28160 46906 28212
rect 2498 28092 2504 28144
rect 2556 28132 2562 28144
rect 2556 28104 44022 28132
rect 2556 28092 2562 28104
rect 45738 28092 45744 28144
rect 45796 28132 45802 28144
rect 46293 28135 46351 28141
rect 46293 28132 46305 28135
rect 45796 28104 46305 28132
rect 45796 28092 45802 28104
rect 46293 28101 46305 28104
rect 46339 28101 46351 28135
rect 46293 28095 46351 28101
rect 54757 28135 54815 28141
rect 54757 28101 54769 28135
rect 54803 28132 54815 28135
rect 57238 28132 57244 28144
rect 54803 28104 57244 28132
rect 54803 28101 54815 28104
rect 54757 28095 54815 28101
rect 57238 28092 57244 28104
rect 57296 28092 57302 28144
rect 44634 28064 44640 28076
rect 44595 28036 44640 28064
rect 44634 28024 44640 28036
rect 44692 28024 44698 28076
rect 45094 28064 45100 28076
rect 45055 28036 45100 28064
rect 45094 28024 45100 28036
rect 45152 28024 45158 28076
rect 45830 28024 45836 28076
rect 45888 28064 45894 28076
rect 46201 28067 46259 28073
rect 46201 28064 46213 28067
rect 45888 28036 46213 28064
rect 45888 28024 45894 28036
rect 46201 28033 46213 28036
rect 46247 28033 46259 28067
rect 46201 28027 46259 28033
rect 46385 28067 46443 28073
rect 46385 28033 46397 28067
rect 46431 28033 46443 28067
rect 47854 28064 47860 28076
rect 47815 28036 47860 28064
rect 46385 28027 46443 28033
rect 46290 27956 46296 28008
rect 46348 27996 46354 28008
rect 46400 27996 46428 28027
rect 47854 28024 47860 28036
rect 47912 28024 47918 28076
rect 47949 28067 48007 28073
rect 47949 28033 47961 28067
rect 47995 28033 48007 28067
rect 48498 28064 48504 28076
rect 48459 28036 48504 28064
rect 47949 28027 48007 28033
rect 46348 27968 46428 27996
rect 46348 27956 46354 27968
rect 47486 27956 47492 28008
rect 47544 27996 47550 28008
rect 47964 27996 47992 28027
rect 48498 28024 48504 28036
rect 48556 28024 48562 28076
rect 49329 28067 49387 28073
rect 49329 28033 49341 28067
rect 49375 28033 49387 28067
rect 49694 28064 49700 28076
rect 49655 28036 49700 28064
rect 49329 28027 49387 28033
rect 47544 27968 47992 27996
rect 48317 27999 48375 28005
rect 47544 27956 47550 27968
rect 48317 27965 48329 27999
rect 48363 27996 48375 27999
rect 49344 27996 49372 28027
rect 49694 28024 49700 28036
rect 49752 28024 49758 28076
rect 50341 28067 50399 28073
rect 50341 28033 50353 28067
rect 50387 28064 50399 28067
rect 50614 28064 50620 28076
rect 50387 28036 50620 28064
rect 50387 28033 50399 28036
rect 50341 28027 50399 28033
rect 50614 28024 50620 28036
rect 50672 28024 50678 28076
rect 50798 28064 50804 28076
rect 50724 28036 50804 28064
rect 49418 27996 49424 28008
rect 48363 27968 49424 27996
rect 48363 27965 48375 27968
rect 48317 27959 48375 27965
rect 49418 27956 49424 27968
rect 49476 27956 49482 28008
rect 49786 27996 49792 28008
rect 49747 27968 49792 27996
rect 49786 27956 49792 27968
rect 49844 27996 49850 28008
rect 50724 27996 50752 28036
rect 50798 28024 50804 28036
rect 50856 28064 50862 28076
rect 51169 28067 51227 28073
rect 51169 28064 51181 28067
rect 50856 28036 51181 28064
rect 50856 28024 50862 28036
rect 51169 28033 51181 28036
rect 51215 28033 51227 28067
rect 51350 28064 51356 28076
rect 51311 28036 51356 28064
rect 51169 28027 51227 28033
rect 51350 28024 51356 28036
rect 51408 28024 51414 28076
rect 52181 28067 52239 28073
rect 52181 28064 52193 28067
rect 51552 28036 52193 28064
rect 51074 27996 51080 28008
rect 49844 27968 50752 27996
rect 51035 27968 51080 27996
rect 49844 27956 49850 27968
rect 51074 27956 51080 27968
rect 51132 27956 51138 28008
rect 51552 28005 51580 28036
rect 52181 28033 52193 28036
rect 52227 28033 52239 28067
rect 52181 28027 52239 28033
rect 52365 28067 52423 28073
rect 52365 28033 52377 28067
rect 52411 28064 52423 28067
rect 52822 28064 52828 28076
rect 52411 28036 52828 28064
rect 52411 28033 52423 28036
rect 52365 28027 52423 28033
rect 52822 28024 52828 28036
rect 52880 28024 52886 28076
rect 52917 28067 52975 28073
rect 52917 28033 52929 28067
rect 52963 28033 52975 28067
rect 52917 28027 52975 28033
rect 51261 27999 51319 28005
rect 51261 27965 51273 27999
rect 51307 27965 51319 27999
rect 51261 27959 51319 27965
rect 51537 27999 51595 28005
rect 51537 27965 51549 27999
rect 51583 27965 51595 27999
rect 52932 27996 52960 28027
rect 53006 28024 53012 28076
rect 53064 28064 53070 28076
rect 53285 28067 53343 28073
rect 53285 28064 53297 28067
rect 53064 28036 53297 28064
rect 53064 28024 53070 28036
rect 53285 28033 53297 28036
rect 53331 28064 53343 28067
rect 53742 28064 53748 28076
rect 53331 28036 53748 28064
rect 53331 28033 53343 28036
rect 53285 28027 53343 28033
rect 53742 28024 53748 28036
rect 53800 28024 53806 28076
rect 54021 28067 54079 28073
rect 54021 28033 54033 28067
rect 54067 28064 54079 28067
rect 54202 28064 54208 28076
rect 54067 28036 54208 28064
rect 54067 28033 54079 28036
rect 54021 28027 54079 28033
rect 54202 28024 54208 28036
rect 54260 28024 54266 28076
rect 54386 28064 54392 28076
rect 54347 28036 54392 28064
rect 54386 28024 54392 28036
rect 54444 28024 54450 28076
rect 54665 28067 54723 28073
rect 54665 28033 54677 28067
rect 54711 28064 54723 28067
rect 55582 28064 55588 28076
rect 54711 28036 55588 28064
rect 54711 28033 54723 28036
rect 54665 28027 54723 28033
rect 55582 28024 55588 28036
rect 55640 28024 55646 28076
rect 55858 28064 55864 28076
rect 55819 28036 55864 28064
rect 55858 28024 55864 28036
rect 55916 28024 55922 28076
rect 56042 28024 56048 28076
rect 56100 28064 56106 28076
rect 56137 28067 56195 28073
rect 56137 28064 56149 28067
rect 56100 28036 56149 28064
rect 56100 28024 56106 28036
rect 56137 28033 56149 28036
rect 56183 28033 56195 28067
rect 56137 28027 56195 28033
rect 53926 27996 53932 28008
rect 52932 27968 53932 27996
rect 51537 27959 51595 27965
rect 45922 27888 45928 27940
rect 45980 27928 45986 27940
rect 46017 27931 46075 27937
rect 46017 27928 46029 27931
rect 45980 27900 46029 27928
rect 45980 27888 45986 27900
rect 46017 27897 46029 27900
rect 46063 27897 46075 27931
rect 46017 27891 46075 27897
rect 50982 27888 50988 27940
rect 51040 27928 51046 27940
rect 51276 27928 51304 27959
rect 53926 27956 53932 27968
rect 53984 27956 53990 28008
rect 55214 27956 55220 28008
rect 55272 27996 55278 28008
rect 55272 27968 55317 27996
rect 55272 27956 55278 27968
rect 51040 27900 51304 27928
rect 51040 27888 51046 27900
rect 47118 27860 47124 27872
rect 47079 27832 47124 27860
rect 47118 27820 47124 27832
rect 47176 27820 47182 27872
rect 52273 27863 52331 27869
rect 52273 27829 52285 27863
rect 52319 27860 52331 27863
rect 53190 27860 53196 27872
rect 52319 27832 53196 27860
rect 52319 27829 52331 27832
rect 52273 27823 52331 27829
rect 53190 27820 53196 27832
rect 53248 27820 53254 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 46014 27616 46020 27668
rect 46072 27656 46078 27668
rect 46109 27659 46167 27665
rect 46109 27656 46121 27659
rect 46072 27628 46121 27656
rect 46072 27616 46078 27628
rect 46109 27625 46121 27628
rect 46155 27625 46167 27659
rect 47210 27656 47216 27668
rect 47171 27628 47216 27656
rect 46109 27619 46167 27625
rect 47210 27616 47216 27628
rect 47268 27616 47274 27668
rect 49237 27659 49295 27665
rect 49237 27625 49249 27659
rect 49283 27656 49295 27659
rect 49602 27656 49608 27668
rect 49283 27628 49608 27656
rect 49283 27625 49295 27628
rect 49237 27619 49295 27625
rect 49602 27616 49608 27628
rect 49660 27616 49666 27668
rect 51077 27659 51135 27665
rect 51077 27625 51089 27659
rect 51123 27656 51135 27659
rect 51350 27656 51356 27668
rect 51123 27628 51356 27656
rect 51123 27625 51135 27628
rect 51077 27619 51135 27625
rect 51350 27616 51356 27628
rect 51408 27616 51414 27668
rect 45646 27588 45652 27600
rect 44008 27560 45652 27588
rect 44008 27464 44036 27560
rect 45646 27548 45652 27560
rect 45704 27548 45710 27600
rect 46845 27591 46903 27597
rect 46845 27557 46857 27591
rect 46891 27588 46903 27591
rect 47854 27588 47860 27600
rect 46891 27560 47860 27588
rect 46891 27557 46903 27560
rect 46845 27551 46903 27557
rect 47854 27548 47860 27560
rect 47912 27548 47918 27600
rect 47946 27548 47952 27600
rect 48004 27588 48010 27600
rect 48225 27591 48283 27597
rect 48225 27588 48237 27591
rect 48004 27560 48237 27588
rect 48004 27548 48010 27560
rect 48225 27557 48237 27560
rect 48271 27557 48283 27591
rect 48225 27551 48283 27557
rect 53745 27591 53803 27597
rect 53745 27557 53757 27591
rect 53791 27588 53803 27591
rect 54202 27588 54208 27600
rect 53791 27560 54208 27588
rect 53791 27557 53803 27560
rect 53745 27551 53803 27557
rect 54202 27548 54208 27560
rect 54260 27548 54266 27600
rect 55582 27588 55588 27600
rect 55543 27560 55588 27588
rect 55582 27548 55588 27560
rect 55640 27548 55646 27600
rect 44634 27520 44640 27532
rect 44595 27492 44640 27520
rect 44634 27480 44640 27492
rect 44692 27480 44698 27532
rect 45922 27520 45928 27532
rect 45572 27492 45928 27520
rect 43898 27452 43904 27464
rect 43859 27424 43904 27452
rect 43898 27412 43904 27424
rect 43956 27412 43962 27464
rect 43990 27412 43996 27464
rect 44048 27452 44054 27464
rect 44174 27452 44180 27464
rect 44048 27424 44093 27452
rect 44135 27424 44180 27452
rect 44048 27412 44054 27424
rect 44174 27412 44180 27424
rect 44232 27412 44238 27464
rect 44450 27412 44456 27464
rect 44508 27452 44514 27464
rect 45572 27452 45600 27492
rect 45922 27480 45928 27492
rect 45980 27480 45986 27532
rect 47486 27480 47492 27532
rect 47544 27520 47550 27532
rect 47765 27523 47823 27529
rect 47765 27520 47777 27523
rect 47544 27492 47777 27520
rect 47544 27480 47550 27492
rect 47765 27489 47777 27492
rect 47811 27489 47823 27523
rect 47765 27483 47823 27489
rect 45738 27452 45744 27464
rect 44508 27424 45600 27452
rect 45699 27424 45744 27452
rect 44508 27412 44514 27424
rect 45738 27412 45744 27424
rect 45796 27412 45802 27464
rect 45830 27412 45836 27464
rect 45888 27452 45894 27464
rect 46109 27455 46167 27461
rect 45888 27424 45933 27452
rect 45888 27412 45894 27424
rect 46109 27421 46121 27455
rect 46155 27452 46167 27455
rect 46290 27452 46296 27464
rect 46155 27424 46296 27452
rect 46155 27421 46167 27424
rect 46109 27415 46167 27421
rect 46290 27412 46296 27424
rect 46348 27412 46354 27464
rect 46658 27412 46664 27464
rect 46716 27452 46722 27464
rect 47029 27455 47087 27461
rect 47029 27452 47041 27455
rect 46716 27424 47041 27452
rect 46716 27412 46722 27424
rect 47029 27421 47041 27424
rect 47075 27421 47087 27455
rect 47029 27415 47087 27421
rect 47213 27455 47271 27461
rect 47213 27421 47225 27455
rect 47259 27452 47271 27455
rect 47302 27452 47308 27464
rect 47259 27424 47308 27452
rect 47259 27421 47271 27424
rect 47213 27415 47271 27421
rect 47302 27412 47308 27424
rect 47360 27412 47366 27464
rect 47872 27461 47900 27548
rect 52270 27520 52276 27532
rect 52231 27492 52276 27520
rect 52270 27480 52276 27492
rect 52328 27480 52334 27532
rect 52914 27520 52920 27532
rect 52875 27492 52920 27520
rect 52914 27480 52920 27492
rect 52972 27480 52978 27532
rect 54386 27520 54392 27532
rect 53668 27492 54392 27520
rect 47857 27455 47915 27461
rect 47857 27421 47869 27455
rect 47903 27421 47915 27455
rect 49418 27452 49424 27464
rect 49379 27424 49424 27452
rect 47857 27415 47915 27421
rect 49418 27412 49424 27424
rect 49476 27412 49482 27464
rect 49694 27452 49700 27464
rect 49655 27424 49700 27452
rect 49694 27412 49700 27424
rect 49752 27412 49758 27464
rect 50614 27452 50620 27464
rect 50575 27424 50620 27452
rect 50614 27412 50620 27424
rect 50672 27412 50678 27464
rect 50890 27452 50896 27464
rect 50851 27424 50896 27452
rect 50890 27412 50896 27424
rect 50948 27412 50954 27464
rect 52362 27452 52368 27464
rect 52323 27424 52368 27452
rect 52362 27412 52368 27424
rect 52420 27412 52426 27464
rect 53668 27461 53696 27492
rect 54386 27480 54392 27492
rect 54444 27480 54450 27532
rect 53653 27455 53711 27461
rect 53653 27421 53665 27455
rect 53699 27421 53711 27455
rect 53653 27415 53711 27421
rect 53742 27412 53748 27464
rect 53800 27452 53806 27464
rect 53837 27455 53895 27461
rect 53837 27452 53849 27455
rect 53800 27424 53849 27452
rect 53800 27412 53806 27424
rect 53837 27421 53849 27424
rect 53883 27421 53895 27455
rect 53837 27415 53895 27421
rect 53926 27412 53932 27464
rect 53984 27452 53990 27464
rect 54110 27452 54116 27464
rect 53984 27424 54029 27452
rect 54071 27424 54116 27452
rect 53984 27412 53990 27424
rect 54110 27412 54116 27424
rect 54168 27412 54174 27464
rect 54570 27452 54576 27464
rect 54531 27424 54576 27452
rect 54570 27412 54576 27424
rect 54628 27412 54634 27464
rect 55214 27412 55220 27464
rect 55272 27452 55278 27464
rect 55493 27455 55551 27461
rect 55493 27452 55505 27455
rect 55272 27424 55505 27452
rect 55272 27412 55278 27424
rect 55493 27421 55505 27424
rect 55539 27421 55551 27455
rect 56962 27452 56968 27464
rect 56923 27424 56968 27452
rect 55493 27415 55551 27421
rect 56962 27412 56968 27424
rect 57020 27412 57026 27464
rect 57882 27452 57888 27464
rect 57843 27424 57888 27452
rect 57882 27412 57888 27424
rect 57940 27412 57946 27464
rect 2406 27344 2412 27396
rect 2464 27384 2470 27396
rect 56413 27387 56471 27393
rect 56413 27384 56425 27387
rect 2464 27356 56425 27384
rect 2464 27344 2470 27356
rect 56413 27353 56425 27356
rect 56459 27353 56471 27387
rect 56413 27347 56471 27353
rect 49510 27276 49516 27328
rect 49568 27316 49574 27328
rect 49605 27319 49663 27325
rect 49605 27316 49617 27319
rect 49568 27288 49617 27316
rect 49568 27276 49574 27288
rect 49605 27285 49617 27288
rect 49651 27285 49663 27319
rect 50706 27316 50712 27328
rect 50667 27288 50712 27316
rect 49605 27279 49663 27285
rect 50706 27276 50712 27288
rect 50764 27276 50770 27328
rect 53926 27276 53932 27328
rect 53984 27316 53990 27328
rect 54665 27319 54723 27325
rect 54665 27316 54677 27319
rect 53984 27288 54677 27316
rect 53984 27276 53990 27288
rect 54665 27285 54677 27288
rect 54711 27285 54723 27319
rect 54665 27279 54723 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 45738 27072 45744 27124
rect 45796 27112 45802 27124
rect 45925 27115 45983 27121
rect 45925 27112 45937 27115
rect 45796 27084 45937 27112
rect 45796 27072 45802 27084
rect 45925 27081 45937 27084
rect 45971 27081 45983 27115
rect 45925 27075 45983 27081
rect 47302 27072 47308 27124
rect 47360 27112 47366 27124
rect 47765 27115 47823 27121
rect 47765 27112 47777 27115
rect 47360 27084 47777 27112
rect 47360 27072 47366 27084
rect 47765 27081 47777 27084
rect 47811 27112 47823 27115
rect 48498 27112 48504 27124
rect 47811 27084 48504 27112
rect 47811 27081 47823 27084
rect 47765 27075 47823 27081
rect 48498 27072 48504 27084
rect 48556 27072 48562 27124
rect 51166 27112 51172 27124
rect 51127 27084 51172 27112
rect 51166 27072 51172 27084
rect 51224 27072 51230 27124
rect 52365 27115 52423 27121
rect 52365 27081 52377 27115
rect 52411 27112 52423 27115
rect 54386 27112 54392 27124
rect 52411 27084 53420 27112
rect 54347 27084 54392 27112
rect 52411 27081 52423 27084
rect 52365 27075 52423 27081
rect 43533 27047 43591 27053
rect 43533 27013 43545 27047
rect 43579 27044 43591 27047
rect 44450 27044 44456 27056
rect 43579 27016 44456 27044
rect 43579 27013 43591 27016
rect 43533 27007 43591 27013
rect 44450 27004 44456 27016
rect 44508 27004 44514 27056
rect 47118 27044 47124 27056
rect 45940 27016 47124 27044
rect 43441 26979 43499 26985
rect 43441 26945 43453 26979
rect 43487 26945 43499 26979
rect 43441 26939 43499 26945
rect 43717 26979 43775 26985
rect 43717 26945 43729 26979
rect 43763 26976 43775 26979
rect 43806 26976 43812 26988
rect 43763 26948 43812 26976
rect 43763 26945 43775 26948
rect 43717 26939 43775 26945
rect 43456 26908 43484 26939
rect 43806 26936 43812 26948
rect 43864 26936 43870 26988
rect 43898 26936 43904 26988
rect 43956 26976 43962 26988
rect 44177 26979 44235 26985
rect 44177 26976 44189 26979
rect 43956 26948 44189 26976
rect 43956 26936 43962 26948
rect 44177 26945 44189 26948
rect 44223 26945 44235 26979
rect 44177 26939 44235 26945
rect 44634 26936 44640 26988
rect 44692 26976 44698 26988
rect 44821 26979 44879 26985
rect 44821 26976 44833 26979
rect 44692 26948 44833 26976
rect 44692 26936 44698 26948
rect 44821 26945 44833 26948
rect 44867 26945 44879 26979
rect 44821 26939 44879 26945
rect 44266 26908 44272 26920
rect 26206 26880 41414 26908
rect 43456 26880 44272 26908
rect 12434 26800 12440 26852
rect 12492 26840 12498 26852
rect 26206 26840 26234 26880
rect 12492 26812 26234 26840
rect 12492 26800 12498 26812
rect 41386 26772 41414 26880
rect 44266 26868 44272 26880
rect 44324 26868 44330 26920
rect 44910 26908 44916 26920
rect 44871 26880 44916 26908
rect 44910 26868 44916 26880
rect 44968 26868 44974 26920
rect 45940 26917 45968 27016
rect 47118 27004 47124 27016
rect 47176 27004 47182 27056
rect 47578 27004 47584 27056
rect 47636 27044 47642 27056
rect 47949 27047 48007 27053
rect 47949 27044 47961 27047
rect 47636 27016 47961 27044
rect 47636 27004 47642 27016
rect 47949 27013 47961 27016
rect 47995 27013 48007 27047
rect 47949 27007 48007 27013
rect 49789 27047 49847 27053
rect 49789 27013 49801 27047
rect 49835 27044 49847 27047
rect 50706 27044 50712 27056
rect 49835 27016 50712 27044
rect 49835 27013 49847 27016
rect 49789 27007 49847 27013
rect 50706 27004 50712 27016
rect 50764 27044 50770 27056
rect 50801 27047 50859 27053
rect 50801 27044 50813 27047
rect 50764 27016 50813 27044
rect 50764 27004 50770 27016
rect 50801 27013 50813 27016
rect 50847 27013 50859 27047
rect 50801 27007 50859 27013
rect 50890 27004 50896 27056
rect 50948 27044 50954 27056
rect 51001 27047 51059 27053
rect 51001 27044 51013 27047
rect 50948 27016 51013 27044
rect 50948 27004 50954 27016
rect 51001 27013 51013 27016
rect 51047 27013 51059 27047
rect 51001 27007 51059 27013
rect 52917 27047 52975 27053
rect 52917 27013 52929 27047
rect 52963 27044 52975 27047
rect 53006 27044 53012 27056
rect 52963 27016 53012 27044
rect 52963 27013 52975 27016
rect 52917 27007 52975 27013
rect 53006 27004 53012 27016
rect 53064 27004 53070 27056
rect 53392 27044 53420 27084
rect 54386 27072 54392 27084
rect 54444 27072 54450 27124
rect 56045 27115 56103 27121
rect 56045 27081 56057 27115
rect 56091 27112 56103 27115
rect 57146 27112 57152 27124
rect 56091 27084 57152 27112
rect 56091 27081 56103 27084
rect 56045 27075 56103 27081
rect 57146 27072 57152 27084
rect 57204 27072 57210 27124
rect 54570 27044 54576 27056
rect 53392 27016 54576 27044
rect 54570 27004 54576 27016
rect 54628 27004 54634 27056
rect 46201 26979 46259 26985
rect 46201 26945 46213 26979
rect 46247 26976 46259 26979
rect 46566 26976 46572 26988
rect 46247 26948 46572 26976
rect 46247 26945 46259 26948
rect 46201 26939 46259 26945
rect 46566 26936 46572 26948
rect 46624 26936 46630 26988
rect 48038 26976 48044 26988
rect 47999 26948 48044 26976
rect 48038 26936 48044 26948
rect 48096 26936 48102 26988
rect 48130 26936 48136 26988
rect 48188 26976 48194 26988
rect 48188 26948 48233 26976
rect 48188 26936 48194 26948
rect 49234 26936 49240 26988
rect 49292 26976 49298 26988
rect 49697 26979 49755 26985
rect 49697 26976 49709 26979
rect 49292 26948 49709 26976
rect 49292 26936 49298 26948
rect 49697 26945 49709 26948
rect 49743 26945 49755 26979
rect 49697 26939 49755 26945
rect 52181 26979 52239 26985
rect 52181 26945 52193 26979
rect 52227 26976 52239 26979
rect 52270 26976 52276 26988
rect 52227 26948 52276 26976
rect 52227 26945 52239 26948
rect 52181 26939 52239 26945
rect 52270 26936 52276 26948
rect 52328 26936 52334 26988
rect 52362 26936 52368 26988
rect 52420 26976 52426 26988
rect 54294 26976 54300 26988
rect 52420 26948 52465 26976
rect 54255 26948 54300 26976
rect 52420 26936 52426 26948
rect 54294 26936 54300 26948
rect 54352 26936 54358 26988
rect 54938 26936 54944 26988
rect 54996 26976 55002 26988
rect 55217 26979 55275 26985
rect 55217 26976 55229 26979
rect 54996 26948 55229 26976
rect 54996 26936 55002 26948
rect 55217 26945 55229 26948
rect 55263 26945 55275 26979
rect 55217 26939 55275 26945
rect 55401 26979 55459 26985
rect 55401 26945 55413 26979
rect 55447 26945 55459 26979
rect 55858 26976 55864 26988
rect 55819 26948 55864 26976
rect 55401 26939 55459 26945
rect 45925 26911 45983 26917
rect 45925 26877 45937 26911
rect 45971 26877 45983 26911
rect 45925 26871 45983 26877
rect 46014 26868 46020 26920
rect 46072 26908 46078 26920
rect 46661 26911 46719 26917
rect 46661 26908 46673 26911
rect 46072 26880 46673 26908
rect 46072 26868 46078 26880
rect 46661 26877 46673 26880
rect 46707 26877 46719 26911
rect 46661 26871 46719 26877
rect 47946 26868 47952 26920
rect 48004 26908 48010 26920
rect 48317 26911 48375 26917
rect 48317 26908 48329 26911
rect 48004 26880 48329 26908
rect 48004 26868 48010 26880
rect 48317 26877 48329 26880
rect 48363 26877 48375 26911
rect 55416 26908 55444 26939
rect 55858 26936 55864 26948
rect 55916 26936 55922 26988
rect 56042 26976 56048 26988
rect 56003 26948 56048 26976
rect 56042 26936 56048 26948
rect 56100 26936 56106 26988
rect 56962 26936 56968 26988
rect 57020 26976 57026 26988
rect 57164 26985 57192 27072
rect 57057 26979 57115 26985
rect 57057 26976 57069 26979
rect 57020 26948 57069 26976
rect 57020 26936 57026 26948
rect 57057 26945 57069 26948
rect 57103 26945 57115 26979
rect 57057 26939 57115 26945
rect 57149 26979 57207 26985
rect 57149 26945 57161 26979
rect 57195 26945 57207 26979
rect 57149 26939 57207 26945
rect 56318 26908 56324 26920
rect 55416 26880 56324 26908
rect 48317 26871 48375 26877
rect 56318 26868 56324 26880
rect 56376 26868 56382 26920
rect 57238 26908 57244 26920
rect 57199 26880 57244 26908
rect 57238 26868 57244 26880
rect 57296 26868 57302 26920
rect 57333 26911 57391 26917
rect 57333 26877 57345 26911
rect 57379 26877 57391 26911
rect 57333 26871 57391 26877
rect 43717 26843 43775 26849
rect 43717 26809 43729 26843
rect 43763 26840 43775 26843
rect 44174 26840 44180 26852
rect 43763 26812 44180 26840
rect 43763 26809 43775 26812
rect 43717 26803 43775 26809
rect 44174 26800 44180 26812
rect 44232 26800 44238 26852
rect 48222 26840 48228 26852
rect 44284 26812 48228 26840
rect 44284 26772 44312 26812
rect 48222 26800 48228 26812
rect 48280 26800 48286 26852
rect 53190 26840 53196 26852
rect 53151 26812 53196 26840
rect 53190 26800 53196 26812
rect 53248 26800 53254 26852
rect 57054 26800 57060 26852
rect 57112 26840 57118 26852
rect 57348 26840 57376 26871
rect 57112 26812 57376 26840
rect 57112 26800 57118 26812
rect 41386 26744 44312 26772
rect 44910 26732 44916 26784
rect 44968 26772 44974 26784
rect 45094 26772 45100 26784
rect 44968 26744 45100 26772
rect 44968 26732 44974 26744
rect 45094 26732 45100 26744
rect 45152 26772 45158 26784
rect 45465 26775 45523 26781
rect 45465 26772 45477 26775
rect 45152 26744 45477 26772
rect 45152 26732 45158 26744
rect 45465 26741 45477 26744
rect 45511 26741 45523 26775
rect 45465 26735 45523 26741
rect 46106 26732 46112 26784
rect 46164 26772 46170 26784
rect 46164 26744 46209 26772
rect 46164 26732 46170 26744
rect 46658 26732 46664 26784
rect 46716 26772 46722 26784
rect 48774 26772 48780 26784
rect 46716 26744 48780 26772
rect 46716 26732 46722 26744
rect 48774 26732 48780 26744
rect 48832 26732 48838 26784
rect 50614 26732 50620 26784
rect 50672 26772 50678 26784
rect 50985 26775 51043 26781
rect 50985 26772 50997 26775
rect 50672 26744 50997 26772
rect 50672 26732 50678 26744
rect 50985 26741 50997 26744
rect 51031 26741 51043 26775
rect 53374 26772 53380 26784
rect 53335 26744 53380 26772
rect 50985 26735 51043 26741
rect 53374 26732 53380 26744
rect 53432 26732 53438 26784
rect 55214 26732 55220 26784
rect 55272 26772 55278 26784
rect 57514 26772 57520 26784
rect 55272 26744 55317 26772
rect 57475 26744 57520 26772
rect 55272 26732 55278 26744
rect 57514 26732 57520 26744
rect 57572 26732 57578 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 43898 26528 43904 26580
rect 43956 26568 43962 26580
rect 44085 26571 44143 26577
rect 44085 26568 44097 26571
rect 43956 26540 44097 26568
rect 43956 26528 43962 26540
rect 44085 26537 44097 26540
rect 44131 26537 44143 26571
rect 44085 26531 44143 26537
rect 44269 26571 44327 26577
rect 44269 26537 44281 26571
rect 44315 26537 44327 26571
rect 44269 26531 44327 26537
rect 45649 26571 45707 26577
rect 45649 26537 45661 26571
rect 45695 26568 45707 26571
rect 46106 26568 46112 26580
rect 45695 26540 46112 26568
rect 45695 26537 45707 26540
rect 45649 26531 45707 26537
rect 38841 26503 38899 26509
rect 38841 26469 38853 26503
rect 38887 26500 38899 26503
rect 40034 26500 40040 26512
rect 38887 26472 40040 26500
rect 38887 26469 38899 26472
rect 38841 26463 38899 26469
rect 40034 26460 40040 26472
rect 40092 26460 40098 26512
rect 43806 26460 43812 26512
rect 43864 26500 43870 26512
rect 44284 26500 44312 26531
rect 46106 26528 46112 26540
rect 46164 26568 46170 26580
rect 46293 26571 46351 26577
rect 46293 26568 46305 26571
rect 46164 26540 46305 26568
rect 46164 26528 46170 26540
rect 46293 26537 46305 26540
rect 46339 26537 46351 26571
rect 47026 26568 47032 26580
rect 46987 26540 47032 26568
rect 46293 26531 46351 26537
rect 47026 26528 47032 26540
rect 47084 26528 47090 26580
rect 47210 26528 47216 26580
rect 47268 26568 47274 26580
rect 47765 26571 47823 26577
rect 47765 26568 47777 26571
rect 47268 26540 47777 26568
rect 47268 26528 47274 26540
rect 47765 26537 47777 26540
rect 47811 26537 47823 26571
rect 47765 26531 47823 26537
rect 49605 26571 49663 26577
rect 49605 26537 49617 26571
rect 49651 26568 49663 26571
rect 49694 26568 49700 26580
rect 49651 26540 49700 26568
rect 49651 26537 49663 26540
rect 49605 26531 49663 26537
rect 49694 26528 49700 26540
rect 49752 26528 49758 26580
rect 50893 26571 50951 26577
rect 50893 26537 50905 26571
rect 50939 26568 50951 26571
rect 50982 26568 50988 26580
rect 50939 26540 50988 26568
rect 50939 26537 50951 26540
rect 50893 26531 50951 26537
rect 50982 26528 50988 26540
rect 51040 26528 51046 26580
rect 53374 26528 53380 26580
rect 53432 26568 53438 26580
rect 58526 26568 58532 26580
rect 53432 26540 58532 26568
rect 53432 26528 53438 26540
rect 58526 26528 58532 26540
rect 58584 26528 58590 26580
rect 45922 26500 45928 26512
rect 43864 26472 45928 26500
rect 43864 26460 43870 26472
rect 45922 26460 45928 26472
rect 45980 26460 45986 26512
rect 46198 26460 46204 26512
rect 46256 26500 46262 26512
rect 47305 26503 47363 26509
rect 46256 26472 47164 26500
rect 46256 26460 46262 26472
rect 46385 26435 46443 26441
rect 46385 26401 46397 26435
rect 46431 26432 46443 26435
rect 46566 26432 46572 26444
rect 46431 26404 46572 26432
rect 46431 26401 46443 26404
rect 46385 26395 46443 26401
rect 46566 26392 46572 26404
rect 46624 26432 46630 26444
rect 47029 26435 47087 26441
rect 47029 26432 47041 26435
rect 46624 26404 47041 26432
rect 46624 26392 46630 26404
rect 47029 26401 47041 26404
rect 47075 26401 47087 26435
rect 47136 26432 47164 26472
rect 47305 26469 47317 26503
rect 47351 26500 47363 26503
rect 48038 26500 48044 26512
rect 47351 26472 48044 26500
rect 47351 26469 47363 26472
rect 47305 26463 47363 26469
rect 48038 26460 48044 26472
rect 48096 26500 48102 26512
rect 48096 26472 48176 26500
rect 48096 26460 48102 26472
rect 47946 26432 47952 26444
rect 47136 26404 47952 26432
rect 47029 26395 47087 26401
rect 47946 26392 47952 26404
rect 48004 26392 48010 26444
rect 45370 26364 45376 26376
rect 45331 26336 45376 26364
rect 45370 26324 45376 26336
rect 45428 26324 45434 26376
rect 45465 26367 45523 26373
rect 45465 26333 45477 26367
rect 45511 26364 45523 26367
rect 46014 26364 46020 26376
rect 45511 26336 46020 26364
rect 45511 26333 45523 26336
rect 45465 26327 45523 26333
rect 46014 26324 46020 26336
rect 46072 26324 46078 26376
rect 46477 26367 46535 26373
rect 46477 26333 46489 26367
rect 46523 26333 46535 26367
rect 46934 26364 46940 26376
rect 46895 26336 46940 26364
rect 46477 26327 46535 26333
rect 38470 26296 38476 26308
rect 38431 26268 38476 26296
rect 38470 26256 38476 26268
rect 38528 26256 38534 26308
rect 44266 26305 44272 26308
rect 44253 26299 44272 26305
rect 44253 26265 44265 26299
rect 44253 26259 44272 26265
rect 44266 26256 44272 26259
rect 44324 26256 44330 26308
rect 44450 26296 44456 26308
rect 44411 26268 44456 26296
rect 44450 26256 44456 26268
rect 44508 26256 44514 26308
rect 45830 26256 45836 26308
rect 45888 26296 45894 26308
rect 46492 26296 46520 26327
rect 46934 26324 46940 26336
rect 46992 26324 46998 26376
rect 47578 26324 47584 26376
rect 47636 26364 47642 26376
rect 48148 26373 48176 26472
rect 48222 26460 48228 26512
rect 48280 26500 48286 26512
rect 53009 26503 53067 26509
rect 53009 26500 53021 26503
rect 48280 26472 53021 26500
rect 48280 26460 48286 26472
rect 53009 26469 53021 26472
rect 53055 26469 53067 26503
rect 53009 26463 53067 26469
rect 54938 26460 54944 26512
rect 54996 26500 55002 26512
rect 56502 26500 56508 26512
rect 54996 26472 56508 26500
rect 54996 26460 55002 26472
rect 56502 26460 56508 26472
rect 56560 26460 56566 26512
rect 56962 26460 56968 26512
rect 57020 26500 57026 26512
rect 57422 26500 57428 26512
rect 57020 26472 57428 26500
rect 57020 26460 57026 26472
rect 57422 26460 57428 26472
rect 57480 26460 57486 26512
rect 57882 26432 57888 26444
rect 57843 26404 57888 26432
rect 57882 26392 57888 26404
rect 57940 26392 57946 26444
rect 47765 26367 47823 26373
rect 47765 26364 47777 26367
rect 47636 26336 47777 26364
rect 47636 26324 47642 26336
rect 47765 26333 47777 26336
rect 47811 26333 47823 26367
rect 47765 26327 47823 26333
rect 48133 26367 48191 26373
rect 48133 26333 48145 26367
rect 48179 26333 48191 26367
rect 48774 26364 48780 26376
rect 48735 26336 48780 26364
rect 48133 26327 48191 26333
rect 48774 26324 48780 26336
rect 48832 26324 48838 26376
rect 49142 26364 49148 26376
rect 49103 26336 49148 26364
rect 49142 26324 49148 26336
rect 49200 26324 49206 26376
rect 49234 26324 49240 26376
rect 49292 26364 49298 26376
rect 49292 26336 49337 26364
rect 49292 26324 49298 26336
rect 49510 26324 49516 26376
rect 49568 26364 49574 26376
rect 50614 26364 50620 26376
rect 49568 26336 50620 26364
rect 49568 26324 49574 26336
rect 50614 26324 50620 26336
rect 50672 26324 50678 26376
rect 50706 26324 50712 26376
rect 50764 26364 50770 26376
rect 53834 26364 53840 26376
rect 50764 26336 50809 26364
rect 53795 26336 53840 26364
rect 50764 26324 50770 26336
rect 53834 26324 53840 26336
rect 53892 26324 53898 26376
rect 54018 26364 54024 26376
rect 53979 26336 54024 26364
rect 54018 26324 54024 26336
rect 54076 26324 54082 26376
rect 56229 26367 56287 26373
rect 56229 26333 56241 26367
rect 56275 26364 56287 26367
rect 56318 26364 56324 26376
rect 56275 26336 56324 26364
rect 56275 26333 56287 26336
rect 56229 26327 56287 26333
rect 56318 26324 56324 26336
rect 56376 26324 56382 26376
rect 56502 26364 56508 26376
rect 56463 26336 56508 26364
rect 56502 26324 56508 26336
rect 56560 26324 56566 26376
rect 57977 26367 58035 26373
rect 57977 26364 57989 26367
rect 57072 26336 57989 26364
rect 57072 26308 57100 26336
rect 57977 26333 57989 26336
rect 58023 26333 58035 26367
rect 58250 26364 58256 26376
rect 58211 26336 58256 26364
rect 57977 26327 58035 26333
rect 58250 26324 58256 26336
rect 58308 26324 58314 26376
rect 47118 26296 47124 26308
rect 45888 26268 46152 26296
rect 46492 26268 47124 26296
rect 45888 26256 45894 26268
rect 38930 26228 38936 26240
rect 38891 26200 38936 26228
rect 38930 26188 38936 26200
rect 38988 26188 38994 26240
rect 46124 26237 46152 26268
rect 47118 26256 47124 26268
rect 47176 26256 47182 26308
rect 48038 26296 48044 26308
rect 47999 26268 48044 26296
rect 48038 26256 48044 26268
rect 48096 26256 48102 26308
rect 49602 26296 49608 26308
rect 49563 26268 49608 26296
rect 49602 26256 49608 26268
rect 49660 26256 49666 26308
rect 50798 26256 50804 26308
rect 50856 26296 50862 26308
rect 50893 26299 50951 26305
rect 50893 26296 50905 26299
rect 50856 26268 50905 26296
rect 50856 26256 50862 26268
rect 50893 26265 50905 26268
rect 50939 26265 50951 26299
rect 50893 26259 50951 26265
rect 55950 26256 55956 26308
rect 56008 26256 56014 26308
rect 57054 26256 57060 26308
rect 57112 26256 57118 26308
rect 46109 26231 46167 26237
rect 46109 26197 46121 26231
rect 46155 26197 46167 26231
rect 46109 26191 46167 26197
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 44637 26027 44695 26033
rect 44637 25993 44649 26027
rect 44683 26024 44695 26027
rect 44726 26024 44732 26036
rect 44683 25996 44732 26024
rect 44683 25993 44695 25996
rect 44637 25987 44695 25993
rect 44726 25984 44732 25996
rect 44784 25984 44790 26036
rect 46109 26027 46167 26033
rect 46109 25993 46121 26027
rect 46155 26024 46167 26027
rect 46845 26027 46903 26033
rect 46155 25996 46704 26024
rect 46155 25993 46167 25996
rect 46109 25987 46167 25993
rect 44266 25916 44272 25968
rect 44324 25956 44330 25968
rect 45189 25959 45247 25965
rect 45189 25956 45201 25959
rect 44324 25928 45201 25956
rect 44324 25916 44330 25928
rect 45189 25925 45201 25928
rect 45235 25925 45247 25959
rect 45370 25956 45376 25968
rect 45189 25919 45247 25925
rect 45296 25928 45376 25956
rect 38930 25888 38936 25900
rect 38891 25860 38936 25888
rect 38930 25848 38936 25860
rect 38988 25848 38994 25900
rect 39022 25848 39028 25900
rect 39080 25888 39086 25900
rect 43993 25891 44051 25897
rect 39080 25860 39125 25888
rect 39080 25848 39086 25860
rect 43993 25857 44005 25891
rect 44039 25888 44051 25891
rect 44726 25888 44732 25900
rect 44039 25860 44732 25888
rect 44039 25857 44051 25860
rect 43993 25851 44051 25857
rect 44726 25848 44732 25860
rect 44784 25848 44790 25900
rect 45296 25897 45324 25928
rect 45370 25916 45376 25928
rect 45428 25956 45434 25968
rect 45738 25956 45744 25968
rect 45428 25928 45744 25956
rect 45428 25916 45434 25928
rect 45738 25916 45744 25928
rect 45796 25916 45802 25968
rect 45946 25959 46004 25965
rect 45946 25925 45958 25959
rect 45992 25956 46004 25959
rect 45992 25928 46060 25956
rect 45992 25925 46004 25928
rect 45946 25919 46004 25925
rect 45281 25891 45339 25897
rect 45281 25857 45293 25891
rect 45327 25857 45339 25891
rect 45281 25851 45339 25857
rect 43898 25820 43904 25832
rect 43859 25792 43904 25820
rect 43898 25780 43904 25792
rect 43956 25780 43962 25832
rect 46032 25752 46060 25928
rect 46566 25888 46572 25900
rect 46527 25860 46572 25888
rect 46566 25848 46572 25860
rect 46624 25848 46630 25900
rect 46676 25897 46704 25996
rect 46845 25993 46857 26027
rect 46891 26024 46903 26027
rect 48038 26024 48044 26036
rect 46891 25996 48044 26024
rect 46891 25993 46903 25996
rect 46845 25987 46903 25993
rect 48038 25984 48044 25996
rect 48096 25984 48102 26036
rect 54018 26024 54024 26036
rect 53979 25996 54024 26024
rect 54018 25984 54024 25996
rect 54076 25984 54082 26036
rect 57146 25984 57152 26036
rect 57204 25984 57210 26036
rect 48774 25916 48780 25968
rect 48832 25956 48838 25968
rect 49145 25959 49203 25965
rect 49145 25956 49157 25959
rect 48832 25928 49157 25956
rect 48832 25916 48838 25928
rect 49145 25925 49157 25928
rect 49191 25956 49203 25959
rect 49602 25956 49608 25968
rect 49191 25928 49608 25956
rect 49191 25925 49203 25928
rect 49145 25919 49203 25925
rect 49602 25916 49608 25928
rect 49660 25916 49666 25968
rect 57164 25956 57192 25984
rect 57241 25959 57299 25965
rect 57241 25956 57253 25959
rect 57164 25928 57253 25956
rect 57241 25925 57253 25928
rect 57287 25925 57299 25959
rect 58161 25959 58219 25965
rect 58161 25956 58173 25959
rect 57241 25919 57299 25925
rect 57440 25928 58173 25956
rect 57440 25900 57468 25928
rect 58161 25925 58173 25928
rect 58207 25925 58219 25959
rect 58161 25919 58219 25925
rect 46661 25891 46719 25897
rect 46661 25857 46673 25891
rect 46707 25888 46719 25891
rect 46934 25888 46940 25900
rect 46707 25860 46940 25888
rect 46707 25857 46719 25860
rect 46661 25851 46719 25857
rect 46934 25848 46940 25860
rect 46992 25848 46998 25900
rect 48866 25848 48872 25900
rect 48924 25888 48930 25900
rect 49418 25888 49424 25900
rect 48924 25860 49424 25888
rect 48924 25848 48930 25860
rect 49418 25848 49424 25860
rect 49476 25848 49482 25900
rect 49878 25848 49884 25900
rect 49936 25888 49942 25900
rect 50341 25891 50399 25897
rect 50341 25888 50353 25891
rect 49936 25860 50353 25888
rect 49936 25848 49942 25860
rect 50341 25857 50353 25860
rect 50387 25857 50399 25891
rect 50706 25888 50712 25900
rect 50667 25860 50712 25888
rect 50341 25851 50399 25857
rect 50706 25848 50712 25860
rect 50764 25848 50770 25900
rect 50982 25888 50988 25900
rect 50943 25860 50988 25888
rect 50982 25848 50988 25860
rect 51040 25848 51046 25900
rect 52917 25891 52975 25897
rect 52917 25857 52929 25891
rect 52963 25888 52975 25891
rect 53190 25888 53196 25900
rect 52963 25860 53196 25888
rect 52963 25857 52975 25860
rect 52917 25851 52975 25857
rect 53190 25848 53196 25860
rect 53248 25848 53254 25900
rect 54021 25891 54079 25897
rect 54021 25857 54033 25891
rect 54067 25857 54079 25891
rect 54021 25851 54079 25857
rect 54205 25891 54263 25897
rect 54205 25857 54217 25891
rect 54251 25888 54263 25891
rect 54294 25888 54300 25900
rect 54251 25860 54300 25888
rect 54251 25857 54263 25860
rect 54205 25851 54263 25857
rect 46106 25780 46112 25832
rect 46164 25820 46170 25832
rect 46845 25823 46903 25829
rect 46845 25820 46857 25823
rect 46164 25792 46857 25820
rect 46164 25780 46170 25792
rect 46845 25789 46857 25792
rect 46891 25820 46903 25823
rect 47026 25820 47032 25832
rect 46891 25792 47032 25820
rect 46891 25789 46903 25792
rect 46845 25783 46903 25789
rect 47026 25780 47032 25792
rect 47084 25780 47090 25832
rect 49234 25820 49240 25832
rect 49195 25792 49240 25820
rect 49234 25780 49240 25792
rect 49292 25780 49298 25832
rect 50801 25823 50859 25829
rect 50801 25789 50813 25823
rect 50847 25820 50859 25823
rect 52178 25820 52184 25832
rect 50847 25792 52184 25820
rect 50847 25789 50859 25792
rect 50801 25783 50859 25789
rect 52178 25780 52184 25792
rect 52236 25780 52242 25832
rect 52730 25780 52736 25832
rect 52788 25820 52794 25832
rect 53009 25823 53067 25829
rect 53009 25820 53021 25823
rect 52788 25792 53021 25820
rect 52788 25780 52794 25792
rect 53009 25789 53021 25792
rect 53055 25789 53067 25823
rect 54036 25820 54064 25851
rect 54294 25848 54300 25860
rect 54352 25848 54358 25900
rect 54386 25848 54392 25900
rect 54444 25888 54450 25900
rect 54941 25891 54999 25897
rect 54941 25888 54953 25891
rect 54444 25860 54953 25888
rect 54444 25848 54450 25860
rect 54941 25857 54953 25860
rect 54987 25857 54999 25891
rect 54941 25851 54999 25857
rect 55030 25848 55036 25900
rect 55088 25888 55094 25900
rect 56042 25888 56048 25900
rect 55088 25860 55133 25888
rect 56003 25860 56048 25888
rect 55088 25848 55094 25860
rect 56042 25848 56048 25860
rect 56100 25848 56106 25900
rect 57054 25888 57060 25900
rect 57015 25860 57060 25888
rect 57054 25848 57060 25860
rect 57112 25848 57118 25900
rect 57146 25848 57152 25900
rect 57204 25888 57210 25900
rect 57422 25888 57428 25900
rect 57204 25860 57249 25888
rect 57383 25860 57428 25888
rect 57204 25848 57210 25860
rect 57422 25848 57428 25860
rect 57480 25848 57486 25900
rect 57517 25891 57575 25897
rect 57517 25857 57529 25891
rect 57563 25888 57575 25891
rect 57606 25888 57612 25900
rect 57563 25860 57612 25888
rect 57563 25857 57575 25860
rect 57517 25851 57575 25857
rect 57606 25848 57612 25860
rect 57664 25848 57670 25900
rect 58069 25891 58127 25897
rect 58069 25857 58081 25891
rect 58115 25888 58127 25891
rect 58250 25888 58256 25900
rect 58115 25860 58256 25888
rect 58115 25857 58127 25860
rect 58069 25851 58127 25857
rect 54757 25823 54815 25829
rect 54757 25820 54769 25823
rect 54036 25792 54769 25820
rect 53009 25783 53067 25789
rect 54220 25764 54248 25792
rect 54757 25789 54769 25792
rect 54803 25789 54815 25823
rect 54757 25783 54815 25789
rect 55858 25780 55864 25832
rect 55916 25820 55922 25832
rect 56137 25823 56195 25829
rect 56137 25820 56149 25823
rect 55916 25792 56149 25820
rect 55916 25780 55922 25792
rect 56137 25789 56149 25792
rect 56183 25789 56195 25823
rect 58084 25820 58112 25851
rect 58250 25848 58256 25860
rect 58308 25848 58314 25900
rect 56137 25783 56195 25789
rect 56428 25792 58112 25820
rect 47118 25752 47124 25764
rect 46032 25724 47124 25752
rect 47118 25712 47124 25724
rect 47176 25752 47182 25764
rect 47176 25724 47716 25752
rect 47176 25712 47182 25724
rect 47688 25696 47716 25724
rect 49510 25712 49516 25764
rect 49568 25752 49574 25764
rect 49605 25755 49663 25761
rect 49605 25752 49617 25755
rect 49568 25724 49617 25752
rect 49568 25712 49574 25724
rect 49605 25721 49617 25724
rect 49651 25721 49663 25755
rect 49605 25715 49663 25721
rect 54202 25712 54208 25764
rect 54260 25712 54266 25764
rect 56428 25761 56456 25792
rect 56413 25755 56471 25761
rect 56413 25721 56425 25755
rect 56459 25721 56471 25755
rect 56413 25715 56471 25721
rect 1946 25644 1952 25696
rect 2004 25684 2010 25696
rect 38105 25687 38163 25693
rect 38105 25684 38117 25687
rect 2004 25656 38117 25684
rect 2004 25644 2010 25656
rect 38105 25653 38117 25656
rect 38151 25653 38163 25687
rect 38105 25647 38163 25653
rect 45925 25687 45983 25693
rect 45925 25653 45937 25687
rect 45971 25684 45983 25687
rect 46014 25684 46020 25696
rect 45971 25656 46020 25684
rect 45971 25653 45983 25656
rect 45925 25647 45983 25653
rect 46014 25644 46020 25656
rect 46072 25644 46078 25696
rect 47670 25644 47676 25696
rect 47728 25684 47734 25696
rect 47765 25687 47823 25693
rect 47765 25684 47777 25687
rect 47728 25656 47777 25684
rect 47728 25644 47734 25656
rect 47765 25653 47777 25656
rect 47811 25684 47823 25687
rect 48317 25687 48375 25693
rect 48317 25684 48329 25687
rect 47811 25656 48329 25684
rect 47811 25653 47823 25656
rect 47765 25647 47823 25653
rect 48317 25653 48329 25656
rect 48363 25653 48375 25687
rect 49142 25684 49148 25696
rect 49103 25656 49148 25684
rect 48317 25647 48375 25653
rect 49142 25644 49148 25656
rect 49200 25644 49206 25696
rect 52454 25644 52460 25696
rect 52512 25684 52518 25696
rect 52917 25687 52975 25693
rect 52917 25684 52929 25687
rect 52512 25656 52929 25684
rect 52512 25644 52518 25656
rect 52917 25653 52929 25656
rect 52963 25653 52975 25687
rect 53282 25684 53288 25696
rect 53243 25656 53288 25684
rect 52917 25647 52975 25653
rect 53282 25644 53288 25656
rect 53340 25644 53346 25696
rect 55214 25644 55220 25696
rect 55272 25684 55278 25696
rect 55950 25684 55956 25696
rect 55272 25656 55956 25684
rect 55272 25644 55278 25656
rect 55950 25644 55956 25656
rect 56008 25684 56014 25696
rect 56045 25687 56103 25693
rect 56045 25684 56057 25687
rect 56008 25656 56057 25684
rect 56008 25644 56014 25656
rect 56045 25653 56057 25656
rect 56091 25653 56103 25687
rect 56870 25684 56876 25696
rect 56831 25656 56876 25684
rect 56045 25647 56103 25653
rect 56870 25644 56876 25656
rect 56928 25644 56934 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 40402 25480 40408 25492
rect 40363 25452 40408 25480
rect 40402 25440 40408 25452
rect 40460 25440 40466 25492
rect 43898 25480 43904 25492
rect 43859 25452 43904 25480
rect 43898 25440 43904 25452
rect 43956 25440 43962 25492
rect 45186 25440 45192 25492
rect 45244 25480 45250 25492
rect 45465 25483 45523 25489
rect 45465 25480 45477 25483
rect 45244 25452 45477 25480
rect 45244 25440 45250 25452
rect 45465 25449 45477 25452
rect 45511 25449 45523 25483
rect 45465 25443 45523 25449
rect 46014 25440 46020 25492
rect 46072 25480 46078 25492
rect 46201 25483 46259 25489
rect 46201 25480 46213 25483
rect 46072 25452 46213 25480
rect 46072 25440 46078 25452
rect 46201 25449 46213 25452
rect 46247 25449 46259 25483
rect 47486 25480 47492 25492
rect 47447 25452 47492 25480
rect 46201 25443 46259 25449
rect 47486 25440 47492 25452
rect 47544 25440 47550 25492
rect 48774 25480 48780 25492
rect 48735 25452 48780 25480
rect 48774 25440 48780 25452
rect 48832 25440 48838 25492
rect 50798 25480 50804 25492
rect 50759 25452 50804 25480
rect 50798 25440 50804 25452
rect 50856 25440 50862 25492
rect 53929 25483 53987 25489
rect 53929 25449 53941 25483
rect 53975 25480 53987 25483
rect 54294 25480 54300 25492
rect 53975 25452 54300 25480
rect 53975 25449 53987 25452
rect 53929 25443 53987 25449
rect 54294 25440 54300 25452
rect 54352 25440 54358 25492
rect 55950 25480 55956 25492
rect 55911 25452 55956 25480
rect 55950 25440 55956 25452
rect 56008 25440 56014 25492
rect 56045 25483 56103 25489
rect 56045 25449 56057 25483
rect 56091 25480 56103 25483
rect 57054 25480 57060 25492
rect 56091 25452 57060 25480
rect 56091 25449 56103 25452
rect 56045 25443 56103 25449
rect 57054 25440 57060 25452
rect 57112 25440 57118 25492
rect 57790 25480 57796 25492
rect 57164 25452 57796 25480
rect 38933 25415 38991 25421
rect 38933 25381 38945 25415
rect 38979 25412 38991 25415
rect 57164 25412 57192 25452
rect 57790 25440 57796 25452
rect 57848 25440 57854 25492
rect 38979 25384 57192 25412
rect 38979 25381 38991 25384
rect 38933 25375 38991 25381
rect 57606 25372 57612 25424
rect 57664 25372 57670 25424
rect 37257 25347 37315 25353
rect 37257 25313 37269 25347
rect 37303 25344 37315 25347
rect 38381 25347 38439 25353
rect 37303 25316 38056 25344
rect 37303 25313 37315 25316
rect 37257 25307 37315 25313
rect 38028 25288 38056 25316
rect 38381 25313 38393 25347
rect 38427 25344 38439 25347
rect 39022 25344 39028 25356
rect 38427 25316 39028 25344
rect 38427 25313 38439 25316
rect 38381 25307 38439 25313
rect 39022 25304 39028 25316
rect 39080 25304 39086 25356
rect 44450 25304 44456 25356
rect 44508 25344 44514 25356
rect 45373 25347 45431 25353
rect 45373 25344 45385 25347
rect 44508 25316 45385 25344
rect 44508 25304 44514 25316
rect 45373 25313 45385 25316
rect 45419 25344 45431 25347
rect 46198 25344 46204 25356
rect 45419 25316 46204 25344
rect 45419 25313 45431 25316
rect 45373 25307 45431 25313
rect 46198 25304 46204 25316
rect 46256 25304 46262 25356
rect 47302 25344 47308 25356
rect 47263 25316 47308 25344
rect 47302 25304 47308 25316
rect 47360 25304 47366 25356
rect 48593 25347 48651 25353
rect 48593 25313 48605 25347
rect 48639 25344 48651 25347
rect 49329 25347 49387 25353
rect 49329 25344 49341 25347
rect 48639 25316 49341 25344
rect 48639 25313 48651 25316
rect 48593 25307 48651 25313
rect 49329 25313 49341 25316
rect 49375 25313 49387 25347
rect 49329 25307 49387 25313
rect 50617 25347 50675 25353
rect 50617 25313 50629 25347
rect 50663 25344 50675 25347
rect 50706 25344 50712 25356
rect 50663 25316 50712 25344
rect 50663 25313 50675 25316
rect 50617 25307 50675 25313
rect 50706 25304 50712 25316
rect 50764 25304 50770 25356
rect 52181 25347 52239 25353
rect 52181 25313 52193 25347
rect 52227 25344 52239 25347
rect 52362 25344 52368 25356
rect 52227 25316 52368 25344
rect 52227 25313 52239 25316
rect 52181 25307 52239 25313
rect 52362 25304 52368 25316
rect 52420 25304 52426 25356
rect 52822 25344 52828 25356
rect 52783 25316 52828 25344
rect 52822 25304 52828 25316
rect 52880 25304 52886 25356
rect 54386 25344 54392 25356
rect 53944 25316 54392 25344
rect 53944 25288 53972 25316
rect 54386 25304 54392 25316
rect 54444 25304 54450 25356
rect 56134 25344 56140 25356
rect 56095 25316 56140 25344
rect 56134 25304 56140 25316
rect 56192 25304 56198 25356
rect 57624 25344 57652 25372
rect 58069 25347 58127 25353
rect 58069 25344 58081 25347
rect 57624 25316 58081 25344
rect 58069 25313 58081 25316
rect 58115 25313 58127 25347
rect 58069 25307 58127 25313
rect 37461 25279 37519 25285
rect 37461 25245 37473 25279
rect 37507 25276 37519 25279
rect 37734 25276 37740 25288
rect 37507 25248 37740 25276
rect 37507 25245 37519 25248
rect 37461 25239 37519 25245
rect 37734 25236 37740 25248
rect 37792 25236 37798 25288
rect 38010 25276 38016 25288
rect 37971 25248 38016 25276
rect 38010 25236 38016 25248
rect 38068 25236 38074 25288
rect 38194 25276 38200 25288
rect 38155 25248 38200 25276
rect 38194 25236 38200 25248
rect 38252 25236 38258 25288
rect 38838 25276 38844 25288
rect 38799 25248 38844 25276
rect 38838 25236 38844 25248
rect 38896 25236 38902 25288
rect 39206 25276 39212 25288
rect 39167 25248 39212 25276
rect 39206 25236 39212 25248
rect 39264 25236 39270 25288
rect 39390 25276 39396 25288
rect 39351 25248 39396 25276
rect 39390 25236 39396 25248
rect 39448 25236 39454 25288
rect 40034 25276 40040 25288
rect 39995 25248 40040 25276
rect 40034 25236 40040 25248
rect 40092 25236 40098 25288
rect 40218 25276 40224 25288
rect 40179 25248 40224 25276
rect 40218 25236 40224 25248
rect 40276 25236 40282 25288
rect 43717 25279 43775 25285
rect 43717 25245 43729 25279
rect 43763 25245 43775 25279
rect 43717 25239 43775 25245
rect 43901 25279 43959 25285
rect 43901 25245 43913 25279
rect 43947 25276 43959 25279
rect 44910 25276 44916 25288
rect 43947 25248 44916 25276
rect 43947 25245 43959 25248
rect 43901 25239 43959 25245
rect 37182 25208 37188 25220
rect 37143 25180 37188 25208
rect 37182 25168 37188 25180
rect 37240 25168 37246 25220
rect 43732 25208 43760 25239
rect 44910 25236 44916 25248
rect 44968 25236 44974 25288
rect 45741 25279 45799 25285
rect 45741 25245 45753 25279
rect 45787 25276 45799 25279
rect 45830 25276 45836 25288
rect 45787 25248 45836 25276
rect 45787 25245 45799 25248
rect 45741 25239 45799 25245
rect 45830 25236 45836 25248
rect 45888 25236 45894 25288
rect 47213 25279 47271 25285
rect 47213 25245 47225 25279
rect 47259 25245 47271 25279
rect 48498 25276 48504 25288
rect 48459 25248 48504 25276
rect 47213 25239 47271 25245
rect 47118 25208 47124 25220
rect 43732 25180 44128 25208
rect 44100 25152 44128 25180
rect 44376 25180 47124 25208
rect 37369 25143 37427 25149
rect 37369 25109 37381 25143
rect 37415 25140 37427 25143
rect 37458 25140 37464 25152
rect 37415 25112 37464 25140
rect 37415 25109 37427 25112
rect 37369 25103 37427 25109
rect 37458 25100 37464 25112
rect 37516 25100 37522 25152
rect 44082 25100 44088 25152
rect 44140 25140 44146 25152
rect 44376 25149 44404 25180
rect 47118 25168 47124 25180
rect 47176 25168 47182 25220
rect 44361 25143 44419 25149
rect 44361 25140 44373 25143
rect 44140 25112 44373 25140
rect 44140 25100 44146 25112
rect 44361 25109 44373 25112
rect 44407 25109 44419 25143
rect 44361 25103 44419 25109
rect 45462 25100 45468 25152
rect 45520 25140 45526 25152
rect 45557 25143 45615 25149
rect 45557 25140 45569 25143
rect 45520 25112 45569 25140
rect 45520 25100 45526 25112
rect 45557 25109 45569 25112
rect 45603 25109 45615 25143
rect 45557 25103 45615 25109
rect 45646 25100 45652 25152
rect 45704 25140 45710 25152
rect 47228 25140 47256 25239
rect 48498 25236 48504 25248
rect 48556 25236 48562 25288
rect 49510 25276 49516 25288
rect 49471 25248 49516 25276
rect 49510 25236 49516 25248
rect 49568 25236 49574 25288
rect 49789 25279 49847 25285
rect 49789 25245 49801 25279
rect 49835 25245 49847 25279
rect 49789 25239 49847 25245
rect 50525 25279 50583 25285
rect 50525 25245 50537 25279
rect 50571 25276 50583 25279
rect 50982 25276 50988 25288
rect 50571 25248 50988 25276
rect 50571 25245 50583 25248
rect 50525 25239 50583 25245
rect 48958 25168 48964 25220
rect 49016 25208 49022 25220
rect 49804 25208 49832 25239
rect 50982 25236 50988 25248
rect 51040 25236 51046 25288
rect 52917 25279 52975 25285
rect 52917 25245 52929 25279
rect 52963 25276 52975 25279
rect 53282 25276 53288 25288
rect 52963 25248 53288 25276
rect 52963 25245 52975 25248
rect 52917 25239 52975 25245
rect 53282 25236 53288 25248
rect 53340 25236 53346 25288
rect 53926 25276 53932 25288
rect 53839 25248 53932 25276
rect 53926 25236 53932 25248
rect 53984 25236 53990 25288
rect 54113 25279 54171 25285
rect 54113 25245 54125 25279
rect 54159 25276 54171 25279
rect 54202 25276 54208 25288
rect 54159 25248 54208 25276
rect 54159 25245 54171 25248
rect 54113 25239 54171 25245
rect 54202 25236 54208 25248
rect 54260 25276 54266 25288
rect 55030 25276 55036 25288
rect 54260 25248 55036 25276
rect 54260 25236 54266 25248
rect 55030 25236 55036 25248
rect 55088 25236 55094 25288
rect 55858 25276 55864 25288
rect 55819 25248 55864 25276
rect 55858 25236 55864 25248
rect 55916 25236 55922 25288
rect 57514 25236 57520 25288
rect 57572 25276 57578 25288
rect 57572 25248 57638 25276
rect 57572 25236 57578 25248
rect 49016 25180 49832 25208
rect 49016 25168 49022 25180
rect 57054 25168 57060 25220
rect 57112 25208 57118 25220
rect 57241 25211 57299 25217
rect 57241 25208 57253 25211
rect 57112 25180 57253 25208
rect 57112 25168 57118 25180
rect 57241 25177 57253 25180
rect 57287 25177 57299 25211
rect 57241 25171 57299 25177
rect 49697 25143 49755 25149
rect 49697 25140 49709 25143
rect 45704 25112 45749 25140
rect 47228 25112 49709 25140
rect 45704 25100 45710 25112
rect 49697 25109 49709 25112
rect 49743 25140 49755 25143
rect 49786 25140 49792 25152
rect 49743 25112 49792 25140
rect 49743 25109 49755 25112
rect 49697 25103 49755 25109
rect 49786 25100 49792 25112
rect 49844 25100 49850 25152
rect 56781 25143 56839 25149
rect 56781 25109 56793 25143
rect 56827 25140 56839 25143
rect 58434 25140 58440 25152
rect 56827 25112 58440 25140
rect 56827 25109 56839 25112
rect 56781 25103 56839 25109
rect 58434 25100 58440 25112
rect 58492 25100 58498 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 36449 24939 36507 24945
rect 36449 24905 36461 24939
rect 36495 24936 36507 24939
rect 37182 24936 37188 24948
rect 36495 24908 37188 24936
rect 36495 24905 36507 24908
rect 36449 24899 36507 24905
rect 37182 24896 37188 24908
rect 37240 24936 37246 24948
rect 37661 24939 37719 24945
rect 37661 24936 37673 24939
rect 37240 24908 37673 24936
rect 37240 24896 37246 24908
rect 37661 24905 37673 24908
rect 37707 24905 37719 24939
rect 37661 24899 37719 24905
rect 37829 24939 37887 24945
rect 37829 24905 37841 24939
rect 37875 24936 37887 24939
rect 38194 24936 38200 24948
rect 37875 24908 38200 24936
rect 37875 24905 37887 24908
rect 37829 24899 37887 24905
rect 38194 24896 38200 24908
rect 38252 24896 38258 24948
rect 38749 24939 38807 24945
rect 38749 24905 38761 24939
rect 38795 24936 38807 24939
rect 40218 24936 40224 24948
rect 38795 24908 39068 24936
rect 40179 24908 40224 24936
rect 38795 24905 38807 24908
rect 38749 24899 38807 24905
rect 37458 24868 37464 24880
rect 37419 24840 37464 24868
rect 37458 24828 37464 24840
rect 37516 24828 37522 24880
rect 38212 24868 38240 24896
rect 38212 24840 38884 24868
rect 35161 24803 35219 24809
rect 35161 24769 35173 24803
rect 35207 24800 35219 24803
rect 35342 24800 35348 24812
rect 35207 24772 35348 24800
rect 35207 24769 35219 24772
rect 35161 24763 35219 24769
rect 35342 24760 35348 24772
rect 35400 24760 35406 24812
rect 36081 24803 36139 24809
rect 36081 24769 36093 24803
rect 36127 24800 36139 24803
rect 36446 24800 36452 24812
rect 36127 24772 36452 24800
rect 36127 24769 36139 24772
rect 36081 24763 36139 24769
rect 36446 24760 36452 24772
rect 36504 24760 36510 24812
rect 38378 24760 38384 24812
rect 38436 24800 38442 24812
rect 38657 24803 38715 24809
rect 38657 24800 38669 24803
rect 38436 24772 38669 24800
rect 38436 24760 38442 24772
rect 38657 24769 38669 24772
rect 38703 24769 38715 24803
rect 38856 24800 38884 24840
rect 38933 24803 38991 24809
rect 38933 24800 38945 24803
rect 38856 24772 38945 24800
rect 38657 24763 38715 24769
rect 38933 24769 38945 24772
rect 38979 24769 38991 24803
rect 39040 24800 39068 24908
rect 40218 24896 40224 24908
rect 40276 24896 40282 24948
rect 47302 24896 47308 24948
rect 47360 24936 47366 24948
rect 47765 24939 47823 24945
rect 47765 24936 47777 24939
rect 47360 24908 47777 24936
rect 47360 24896 47366 24908
rect 47765 24905 47777 24908
rect 47811 24905 47823 24939
rect 47765 24899 47823 24905
rect 48498 24896 48504 24948
rect 48556 24936 48562 24948
rect 48977 24939 49035 24945
rect 48977 24936 48989 24939
rect 48556 24908 48989 24936
rect 48556 24896 48562 24908
rect 48977 24905 48989 24908
rect 49023 24905 49035 24939
rect 48977 24899 49035 24905
rect 49418 24896 49424 24948
rect 49476 24936 49482 24948
rect 50525 24939 50583 24945
rect 49476 24908 50200 24936
rect 49476 24896 49482 24908
rect 44637 24871 44695 24877
rect 44637 24837 44649 24871
rect 44683 24868 44695 24871
rect 44910 24868 44916 24880
rect 44683 24840 44916 24868
rect 44683 24837 44695 24840
rect 44637 24831 44695 24837
rect 44910 24828 44916 24840
rect 44968 24828 44974 24880
rect 46385 24871 46443 24877
rect 46385 24868 46397 24871
rect 45664 24840 46397 24868
rect 39040 24772 39436 24800
rect 38933 24763 38991 24769
rect 31662 24692 31668 24744
rect 31720 24732 31726 24744
rect 34790 24732 34796 24744
rect 31720 24704 34796 24732
rect 31720 24692 31726 24704
rect 34790 24692 34796 24704
rect 34848 24732 34854 24744
rect 34885 24735 34943 24741
rect 34885 24732 34897 24735
rect 34848 24704 34897 24732
rect 34848 24692 34854 24704
rect 34885 24701 34897 24704
rect 34931 24701 34943 24735
rect 34885 24695 34943 24701
rect 36173 24735 36231 24741
rect 36173 24701 36185 24735
rect 36219 24732 36231 24735
rect 36354 24732 36360 24744
rect 36219 24704 36360 24732
rect 36219 24701 36231 24704
rect 36173 24695 36231 24701
rect 36354 24692 36360 24704
rect 36412 24692 36418 24744
rect 39408 24732 39436 24772
rect 39942 24760 39948 24812
rect 40000 24800 40006 24812
rect 40129 24803 40187 24809
rect 40129 24800 40141 24803
rect 40000 24772 40141 24800
rect 40000 24760 40006 24772
rect 40129 24769 40141 24772
rect 40175 24769 40187 24803
rect 40310 24800 40316 24812
rect 40271 24772 40316 24800
rect 40129 24763 40187 24769
rect 40310 24760 40316 24772
rect 40368 24760 40374 24812
rect 43806 24800 43812 24812
rect 43767 24772 43812 24800
rect 43806 24760 43812 24772
rect 43864 24760 43870 24812
rect 45462 24760 45468 24812
rect 45520 24800 45526 24812
rect 45664 24809 45692 24840
rect 46385 24837 46397 24840
rect 46431 24837 46443 24871
rect 46385 24831 46443 24837
rect 47118 24828 47124 24880
rect 47176 24828 47182 24880
rect 48777 24871 48835 24877
rect 47964 24840 48728 24868
rect 45649 24803 45707 24809
rect 45649 24800 45661 24803
rect 45520 24772 45661 24800
rect 45520 24760 45526 24772
rect 45649 24769 45661 24772
rect 45695 24769 45707 24803
rect 45649 24763 45707 24769
rect 45741 24803 45799 24809
rect 45741 24769 45753 24803
rect 45787 24800 45799 24803
rect 46198 24800 46204 24812
rect 45787 24772 46204 24800
rect 45787 24769 45799 24772
rect 45741 24763 45799 24769
rect 46198 24760 46204 24772
rect 46256 24760 46262 24812
rect 46566 24760 46572 24812
rect 46624 24800 46630 24812
rect 46661 24803 46719 24809
rect 46661 24800 46673 24803
rect 46624 24772 46673 24800
rect 46624 24760 46630 24772
rect 46661 24769 46673 24772
rect 46707 24769 46719 24803
rect 47136 24800 47164 24828
rect 47964 24809 47992 24840
rect 47949 24803 48007 24809
rect 47949 24800 47961 24803
rect 47136 24772 47961 24800
rect 46661 24763 46719 24769
rect 47949 24769 47961 24772
rect 47995 24769 48007 24803
rect 47949 24763 48007 24769
rect 48133 24803 48191 24809
rect 48133 24769 48145 24803
rect 48179 24769 48191 24803
rect 48700 24800 48728 24840
rect 48777 24837 48789 24871
rect 48823 24868 48835 24871
rect 49786 24868 49792 24880
rect 48823 24840 49792 24868
rect 48823 24837 48835 24840
rect 48777 24831 48835 24837
rect 49786 24828 49792 24840
rect 49844 24828 49850 24880
rect 50172 24868 50200 24908
rect 50525 24905 50537 24939
rect 50571 24936 50583 24939
rect 50982 24936 50988 24948
rect 50571 24908 50988 24936
rect 50571 24905 50583 24908
rect 50525 24899 50583 24905
rect 50982 24896 50988 24908
rect 51040 24896 51046 24948
rect 52730 24868 52736 24880
rect 50172 24840 50292 24868
rect 49510 24800 49516 24812
rect 48700 24772 49516 24800
rect 48133 24763 48191 24769
rect 40034 24732 40040 24744
rect 39408 24704 40040 24732
rect 40034 24692 40040 24704
rect 40092 24692 40098 24744
rect 45554 24732 45560 24744
rect 45515 24704 45560 24732
rect 45554 24692 45560 24704
rect 45612 24692 45618 24744
rect 45830 24692 45836 24744
rect 45888 24732 45894 24744
rect 45888 24704 45933 24732
rect 45888 24692 45894 24704
rect 46014 24692 46020 24744
rect 46072 24732 46078 24744
rect 46385 24735 46443 24741
rect 46385 24732 46397 24735
rect 46072 24704 46397 24732
rect 46072 24692 46078 24704
rect 46385 24701 46397 24704
rect 46431 24732 46443 24735
rect 47121 24735 47179 24741
rect 47121 24732 47133 24735
rect 46431 24704 47133 24732
rect 46431 24701 46443 24704
rect 46385 24695 46443 24701
rect 47121 24701 47133 24704
rect 47167 24701 47179 24735
rect 47121 24695 47179 24701
rect 34977 24667 35035 24673
rect 34977 24633 34989 24667
rect 35023 24664 35035 24667
rect 35618 24664 35624 24676
rect 35023 24636 35624 24664
rect 35023 24633 35035 24636
rect 34977 24627 35035 24633
rect 35618 24624 35624 24636
rect 35676 24624 35682 24676
rect 38838 24664 38844 24676
rect 37108 24636 38844 24664
rect 35345 24599 35403 24605
rect 35345 24565 35357 24599
rect 35391 24596 35403 24599
rect 37108 24596 37136 24636
rect 38838 24624 38844 24636
rect 38896 24624 38902 24676
rect 38933 24667 38991 24673
rect 38933 24633 38945 24667
rect 38979 24664 38991 24667
rect 39390 24664 39396 24676
rect 38979 24636 39396 24664
rect 38979 24633 38991 24636
rect 38933 24627 38991 24633
rect 39390 24624 39396 24636
rect 39448 24624 39454 24676
rect 44266 24664 44272 24676
rect 44227 24636 44272 24664
rect 44266 24624 44272 24636
rect 44324 24624 44330 24676
rect 44821 24667 44879 24673
rect 44821 24633 44833 24667
rect 44867 24664 44879 24667
rect 48148 24664 48176 24763
rect 49510 24760 49516 24772
rect 49568 24800 49574 24812
rect 49697 24803 49755 24809
rect 49697 24800 49709 24803
rect 49568 24772 49709 24800
rect 49568 24760 49574 24772
rect 49697 24769 49709 24772
rect 49743 24769 49755 24803
rect 49697 24763 49755 24769
rect 49712 24732 49740 24763
rect 49878 24760 49884 24812
rect 49936 24800 49942 24812
rect 50264 24809 50292 24840
rect 52196 24840 52736 24868
rect 52196 24809 52224 24840
rect 52730 24828 52736 24840
rect 52788 24828 52794 24880
rect 50157 24803 50215 24809
rect 50157 24800 50169 24803
rect 49936 24772 50169 24800
rect 49936 24760 49942 24772
rect 50157 24769 50169 24772
rect 50203 24769 50215 24803
rect 50157 24763 50215 24769
rect 50249 24803 50307 24809
rect 50249 24769 50261 24803
rect 50295 24800 50307 24803
rect 52181 24803 52239 24809
rect 52181 24800 52193 24803
rect 50295 24772 52193 24800
rect 50295 24769 50307 24772
rect 50249 24763 50307 24769
rect 52181 24769 52193 24772
rect 52227 24769 52239 24803
rect 52181 24763 52239 24769
rect 52365 24803 52423 24809
rect 52365 24769 52377 24803
rect 52411 24800 52423 24803
rect 52454 24800 52460 24812
rect 52411 24772 52460 24800
rect 52411 24769 52423 24772
rect 52365 24763 52423 24769
rect 52454 24760 52460 24772
rect 52512 24760 52518 24812
rect 52914 24800 52920 24812
rect 52875 24772 52920 24800
rect 52914 24760 52920 24772
rect 52972 24760 52978 24812
rect 53009 24803 53067 24809
rect 53009 24769 53021 24803
rect 53055 24769 53067 24803
rect 53190 24800 53196 24812
rect 53151 24772 53196 24800
rect 53009 24763 53067 24769
rect 49970 24732 49976 24744
rect 49712 24704 49976 24732
rect 49970 24692 49976 24704
rect 50028 24692 50034 24744
rect 52273 24735 52331 24741
rect 52273 24701 52285 24735
rect 52319 24732 52331 24735
rect 53024 24732 53052 24763
rect 53190 24760 53196 24772
rect 53248 24760 53254 24812
rect 53377 24803 53435 24809
rect 53377 24769 53389 24803
rect 53423 24800 53435 24803
rect 53926 24800 53932 24812
rect 53423 24772 53932 24800
rect 53423 24769 53435 24772
rect 53377 24763 53435 24769
rect 53926 24760 53932 24772
rect 53984 24760 53990 24812
rect 54754 24800 54760 24812
rect 54715 24772 54760 24800
rect 54754 24760 54760 24772
rect 54812 24760 54818 24812
rect 55490 24800 55496 24812
rect 55451 24772 55496 24800
rect 55490 24760 55496 24772
rect 55548 24760 55554 24812
rect 56318 24760 56324 24812
rect 56376 24800 56382 24812
rect 57057 24803 57115 24809
rect 57057 24800 57069 24803
rect 56376 24772 57069 24800
rect 56376 24760 56382 24772
rect 57057 24769 57069 24772
rect 57103 24769 57115 24803
rect 57057 24763 57115 24769
rect 57241 24803 57299 24809
rect 57241 24769 57253 24803
rect 57287 24769 57299 24803
rect 57241 24763 57299 24769
rect 58069 24803 58127 24809
rect 58069 24769 58081 24803
rect 58115 24800 58127 24803
rect 58434 24800 58440 24812
rect 58115 24772 58440 24800
rect 58115 24769 58127 24772
rect 58069 24763 58127 24769
rect 56410 24732 56416 24744
rect 52319 24704 53052 24732
rect 56371 24704 56416 24732
rect 52319 24701 52331 24704
rect 52273 24695 52331 24701
rect 56410 24692 56416 24704
rect 56468 24692 56474 24744
rect 56502 24692 56508 24744
rect 56560 24732 56566 24744
rect 57256 24732 57284 24763
rect 58434 24760 58440 24772
rect 58492 24760 58498 24812
rect 56560 24704 57284 24732
rect 56560 24692 56566 24704
rect 44867 24636 48176 24664
rect 44867 24633 44879 24636
rect 44821 24627 44879 24633
rect 35391 24568 37136 24596
rect 37645 24599 37703 24605
rect 35391 24565 35403 24568
rect 35345 24559 35403 24565
rect 37645 24565 37657 24599
rect 37691 24596 37703 24599
rect 37734 24596 37740 24608
rect 37691 24568 37740 24596
rect 37691 24565 37703 24568
rect 37645 24559 37703 24565
rect 37734 24556 37740 24568
rect 37792 24556 37798 24608
rect 43809 24599 43867 24605
rect 43809 24565 43821 24599
rect 43855 24596 43867 24599
rect 43898 24596 43904 24608
rect 43855 24568 43904 24596
rect 43855 24565 43867 24568
rect 43809 24559 43867 24565
rect 43898 24556 43904 24568
rect 43956 24556 43962 24608
rect 44637 24599 44695 24605
rect 44637 24565 44649 24599
rect 44683 24596 44695 24599
rect 44726 24596 44732 24608
rect 44683 24568 44732 24596
rect 44683 24565 44695 24568
rect 44637 24559 44695 24565
rect 44726 24556 44732 24568
rect 44784 24556 44790 24608
rect 45370 24596 45376 24608
rect 45331 24568 45376 24596
rect 45370 24556 45376 24568
rect 45428 24556 45434 24608
rect 45738 24556 45744 24608
rect 45796 24596 45802 24608
rect 46569 24599 46627 24605
rect 46569 24596 46581 24599
rect 45796 24568 46581 24596
rect 45796 24556 45802 24568
rect 46569 24565 46581 24568
rect 46615 24565 46627 24599
rect 48148 24596 48176 24636
rect 49145 24667 49203 24673
rect 49145 24633 49157 24667
rect 49191 24664 49203 24667
rect 50062 24664 50068 24676
rect 49191 24636 50068 24664
rect 49191 24633 49203 24636
rect 49145 24627 49203 24633
rect 50062 24624 50068 24636
rect 50120 24624 50126 24676
rect 48958 24596 48964 24608
rect 48148 24568 48964 24596
rect 46569 24559 46627 24565
rect 48958 24556 48964 24568
rect 49016 24556 49022 24608
rect 50154 24596 50160 24608
rect 50115 24568 50160 24596
rect 50154 24556 50160 24568
rect 50212 24556 50218 24608
rect 56962 24556 56968 24608
rect 57020 24596 57026 24608
rect 57149 24599 57207 24605
rect 57149 24596 57161 24599
rect 57020 24568 57161 24596
rect 57020 24556 57026 24568
rect 57149 24565 57161 24568
rect 57195 24565 57207 24599
rect 58250 24596 58256 24608
rect 58211 24568 58256 24596
rect 57149 24559 57207 24565
rect 58250 24556 58256 24568
rect 58308 24556 58314 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 35437 24395 35495 24401
rect 35437 24361 35449 24395
rect 35483 24392 35495 24395
rect 35618 24392 35624 24404
rect 35483 24364 35624 24392
rect 35483 24361 35495 24364
rect 35437 24355 35495 24361
rect 35618 24352 35624 24364
rect 35676 24352 35682 24404
rect 36262 24352 36268 24404
rect 36320 24392 36326 24404
rect 36725 24395 36783 24401
rect 36725 24392 36737 24395
rect 36320 24364 36737 24392
rect 36320 24352 36326 24364
rect 36725 24361 36737 24364
rect 36771 24361 36783 24395
rect 36725 24355 36783 24361
rect 37093 24395 37151 24401
rect 37093 24361 37105 24395
rect 37139 24392 37151 24395
rect 37458 24392 37464 24404
rect 37139 24364 37464 24392
rect 37139 24361 37151 24364
rect 37093 24355 37151 24361
rect 37458 24352 37464 24364
rect 37516 24352 37522 24404
rect 38378 24392 38384 24404
rect 38339 24364 38384 24392
rect 38378 24352 38384 24364
rect 38436 24352 38442 24404
rect 40034 24392 40040 24404
rect 39995 24364 40040 24392
rect 40034 24352 40040 24364
rect 40092 24352 40098 24404
rect 43990 24392 43996 24404
rect 43951 24364 43996 24392
rect 43990 24352 43996 24364
rect 44048 24352 44054 24404
rect 45186 24352 45192 24404
rect 45244 24392 45250 24404
rect 45373 24395 45431 24401
rect 45373 24392 45385 24395
rect 45244 24364 45385 24392
rect 45244 24352 45250 24364
rect 45373 24361 45385 24364
rect 45419 24361 45431 24395
rect 45373 24355 45431 24361
rect 47118 24352 47124 24404
rect 47176 24392 47182 24404
rect 47581 24395 47639 24401
rect 47581 24392 47593 24395
rect 47176 24364 47593 24392
rect 47176 24352 47182 24364
rect 47581 24361 47593 24364
rect 47627 24361 47639 24395
rect 47581 24355 47639 24361
rect 50525 24395 50583 24401
rect 50525 24361 50537 24395
rect 50571 24392 50583 24395
rect 50706 24392 50712 24404
rect 50571 24364 50712 24392
rect 50571 24361 50583 24364
rect 50525 24355 50583 24361
rect 50706 24352 50712 24364
rect 50764 24352 50770 24404
rect 55858 24392 55864 24404
rect 55819 24364 55864 24392
rect 55858 24352 55864 24364
rect 55916 24352 55922 24404
rect 57149 24395 57207 24401
rect 57149 24361 57161 24395
rect 57195 24392 57207 24395
rect 58066 24392 58072 24404
rect 57195 24364 58072 24392
rect 57195 24361 57207 24364
rect 57149 24355 57207 24361
rect 58066 24352 58072 24364
rect 58124 24352 58130 24404
rect 43898 24284 43904 24336
rect 43956 24324 43962 24336
rect 53006 24324 53012 24336
rect 43956 24296 53012 24324
rect 43956 24284 43962 24296
rect 34790 24216 34796 24268
rect 34848 24256 34854 24268
rect 35345 24259 35403 24265
rect 35345 24256 35357 24259
rect 34848 24228 35357 24256
rect 34848 24216 34854 24228
rect 35345 24225 35357 24228
rect 35391 24225 35403 24259
rect 35345 24219 35403 24225
rect 38746 24216 38752 24268
rect 38804 24256 38810 24268
rect 40310 24256 40316 24268
rect 38804 24228 40316 24256
rect 38804 24216 38810 24228
rect 40310 24216 40316 24228
rect 40368 24256 40374 24268
rect 43257 24259 43315 24265
rect 40368 24228 40724 24256
rect 40368 24216 40374 24228
rect 27062 24148 27068 24200
rect 27120 24188 27126 24200
rect 27525 24191 27583 24197
rect 27525 24188 27537 24191
rect 27120 24160 27537 24188
rect 27120 24148 27126 24160
rect 27525 24157 27537 24160
rect 27571 24157 27583 24191
rect 27525 24151 27583 24157
rect 27614 24148 27620 24200
rect 27672 24188 27678 24200
rect 27709 24191 27767 24197
rect 27709 24188 27721 24191
rect 27672 24160 27721 24188
rect 27672 24148 27678 24160
rect 27709 24157 27721 24160
rect 27755 24188 27767 24191
rect 31478 24188 31484 24200
rect 27755 24160 31484 24188
rect 27755 24157 27767 24160
rect 27709 24151 27767 24157
rect 31478 24148 31484 24160
rect 31536 24148 31542 24200
rect 31570 24148 31576 24200
rect 31628 24188 31634 24200
rect 31941 24191 31999 24197
rect 31941 24188 31953 24191
rect 31628 24160 31953 24188
rect 31628 24148 31634 24160
rect 31941 24157 31953 24160
rect 31987 24157 31999 24191
rect 32490 24188 32496 24200
rect 32451 24160 32496 24188
rect 31941 24151 31999 24157
rect 32490 24148 32496 24160
rect 32548 24148 32554 24200
rect 35250 24188 35256 24200
rect 35211 24160 35256 24188
rect 35250 24148 35256 24160
rect 35308 24148 35314 24200
rect 36446 24148 36452 24200
rect 36504 24188 36510 24200
rect 36633 24191 36691 24197
rect 36633 24188 36645 24191
rect 36504 24160 36645 24188
rect 36504 24148 36510 24160
rect 36633 24157 36645 24160
rect 36679 24157 36691 24191
rect 36633 24151 36691 24157
rect 38010 24148 38016 24200
rect 38068 24188 38074 24200
rect 38381 24191 38439 24197
rect 38381 24188 38393 24191
rect 38068 24160 38393 24188
rect 38068 24148 38074 24160
rect 38381 24157 38393 24160
rect 38427 24157 38439 24191
rect 38381 24151 38439 24157
rect 38470 24148 38476 24200
rect 38528 24188 38534 24200
rect 38565 24191 38623 24197
rect 38565 24188 38577 24191
rect 38528 24160 38577 24188
rect 38528 24148 38534 24160
rect 38565 24157 38577 24160
rect 38611 24157 38623 24191
rect 38565 24151 38623 24157
rect 40126 24148 40132 24200
rect 40184 24188 40190 24200
rect 40221 24191 40279 24197
rect 40221 24188 40233 24191
rect 40184 24160 40233 24188
rect 40184 24148 40190 24160
rect 40221 24157 40233 24160
rect 40267 24157 40279 24191
rect 40586 24188 40592 24200
rect 40547 24160 40592 24188
rect 40221 24151 40279 24157
rect 40586 24148 40592 24160
rect 40644 24148 40650 24200
rect 40696 24197 40724 24228
rect 43257 24225 43269 24259
rect 43303 24256 43315 24259
rect 43303 24228 43852 24256
rect 43303 24225 43315 24228
rect 43257 24219 43315 24225
rect 43824 24200 43852 24228
rect 40681 24191 40739 24197
rect 40681 24157 40693 24191
rect 40727 24157 40739 24191
rect 40681 24151 40739 24157
rect 43165 24191 43223 24197
rect 43165 24157 43177 24191
rect 43211 24157 43223 24191
rect 43165 24151 43223 24157
rect 43349 24191 43407 24197
rect 43349 24157 43361 24191
rect 43395 24188 43407 24191
rect 43438 24188 43444 24200
rect 43395 24160 43444 24188
rect 43395 24157 43407 24160
rect 43349 24151 43407 24157
rect 10042 24080 10048 24132
rect 10100 24120 10106 24132
rect 40313 24123 40371 24129
rect 40313 24120 40325 24123
rect 10100 24092 32338 24120
rect 40236 24092 40325 24120
rect 10100 24080 10106 24092
rect 40236 24064 40264 24092
rect 40313 24089 40325 24092
rect 40359 24089 40371 24123
rect 40313 24083 40371 24089
rect 40405 24123 40463 24129
rect 40405 24089 40417 24123
rect 40451 24120 40463 24123
rect 41230 24120 41236 24132
rect 40451 24092 41236 24120
rect 40451 24089 40463 24092
rect 40405 24083 40463 24089
rect 41230 24080 41236 24092
rect 41288 24080 41294 24132
rect 43180 24120 43208 24151
rect 43438 24148 43444 24160
rect 43496 24148 43502 24200
rect 43806 24188 43812 24200
rect 43767 24160 43812 24188
rect 43806 24148 43812 24160
rect 43864 24148 43870 24200
rect 44174 24120 44180 24132
rect 43180 24092 44180 24120
rect 44174 24080 44180 24092
rect 44232 24080 44238 24132
rect 45370 24129 45376 24132
rect 45357 24123 45376 24129
rect 45357 24089 45369 24123
rect 45357 24083 45376 24089
rect 45370 24080 45376 24083
rect 45428 24080 45434 24132
rect 45557 24123 45615 24129
rect 45557 24089 45569 24123
rect 45603 24120 45615 24123
rect 45664 24120 45692 24296
rect 53006 24284 53012 24296
rect 53064 24284 53070 24336
rect 50893 24259 50951 24265
rect 50893 24225 50905 24259
rect 50939 24256 50951 24259
rect 51626 24256 51632 24268
rect 50939 24228 51632 24256
rect 50939 24225 50951 24228
rect 50893 24219 50951 24225
rect 51626 24216 51632 24228
rect 51684 24216 51690 24268
rect 54941 24259 54999 24265
rect 54941 24225 54953 24259
rect 54987 24256 54999 24259
rect 55766 24256 55772 24268
rect 54987 24228 55772 24256
rect 54987 24225 54999 24228
rect 54941 24219 54999 24225
rect 55766 24216 55772 24228
rect 55824 24216 55830 24268
rect 56781 24259 56839 24265
rect 56781 24225 56793 24259
rect 56827 24256 56839 24259
rect 57609 24259 57667 24265
rect 57609 24256 57621 24259
rect 56827 24228 57621 24256
rect 56827 24225 56839 24228
rect 56781 24219 56839 24225
rect 57609 24225 57621 24228
rect 57655 24225 57667 24259
rect 57609 24219 57667 24225
rect 46569 24191 46627 24197
rect 46569 24157 46581 24191
rect 46615 24188 46627 24191
rect 46658 24188 46664 24200
rect 46615 24160 46664 24188
rect 46615 24157 46627 24160
rect 46569 24151 46627 24157
rect 46658 24148 46664 24160
rect 46716 24148 46722 24200
rect 46842 24188 46848 24200
rect 46803 24160 46848 24188
rect 46842 24148 46848 24160
rect 46900 24148 46906 24200
rect 50798 24188 50804 24200
rect 50759 24160 50804 24188
rect 50798 24148 50804 24160
rect 50856 24148 50862 24200
rect 52641 24191 52699 24197
rect 52641 24157 52653 24191
rect 52687 24188 52699 24191
rect 52730 24188 52736 24200
rect 52687 24160 52736 24188
rect 52687 24157 52699 24160
rect 52641 24151 52699 24157
rect 52730 24148 52736 24160
rect 52788 24148 52794 24200
rect 53098 24148 53104 24200
rect 53156 24188 53162 24200
rect 53837 24191 53895 24197
rect 53837 24188 53849 24191
rect 53156 24160 53849 24188
rect 53156 24148 53162 24160
rect 53837 24157 53849 24160
rect 53883 24157 53895 24191
rect 53837 24151 53895 24157
rect 53926 24148 53932 24200
rect 53984 24188 53990 24200
rect 54205 24191 54263 24197
rect 54205 24188 54217 24191
rect 53984 24160 54217 24188
rect 53984 24148 53990 24160
rect 54205 24157 54217 24160
rect 54251 24157 54263 24191
rect 54662 24188 54668 24200
rect 54623 24160 54668 24188
rect 54205 24151 54263 24157
rect 54662 24148 54668 24160
rect 54720 24148 54726 24200
rect 55490 24188 55496 24200
rect 55451 24160 55496 24188
rect 55490 24148 55496 24160
rect 55548 24148 55554 24200
rect 55677 24191 55735 24197
rect 55677 24157 55689 24191
rect 55723 24157 55735 24191
rect 55677 24151 55735 24157
rect 45603 24092 45692 24120
rect 46753 24123 46811 24129
rect 45603 24089 45615 24092
rect 45557 24083 45615 24089
rect 46753 24089 46765 24123
rect 46799 24120 46811 24123
rect 46934 24120 46940 24132
rect 46799 24092 46940 24120
rect 46799 24089 46811 24092
rect 46753 24083 46811 24089
rect 46934 24080 46940 24092
rect 46992 24080 46998 24132
rect 52457 24123 52515 24129
rect 52457 24089 52469 24123
rect 52503 24120 52515 24123
rect 52546 24120 52552 24132
rect 52503 24092 52552 24120
rect 52503 24089 52515 24092
rect 52457 24083 52515 24089
rect 52546 24080 52552 24092
rect 52604 24080 52610 24132
rect 54754 24080 54760 24132
rect 54812 24120 54818 24132
rect 55692 24120 55720 24151
rect 56410 24148 56416 24200
rect 56468 24188 56474 24200
rect 56689 24191 56747 24197
rect 56689 24188 56701 24191
rect 56468 24160 56701 24188
rect 56468 24148 56474 24160
rect 56689 24157 56701 24160
rect 56735 24157 56747 24191
rect 56962 24188 56968 24200
rect 56923 24160 56968 24188
rect 56689 24151 56747 24157
rect 56962 24148 56968 24160
rect 57020 24148 57026 24200
rect 57793 24191 57851 24197
rect 57793 24157 57805 24191
rect 57839 24188 57851 24191
rect 57882 24188 57888 24200
rect 57839 24160 57888 24188
rect 57839 24157 57851 24160
rect 57793 24151 57851 24157
rect 57882 24148 57888 24160
rect 57940 24148 57946 24200
rect 58066 24188 58072 24200
rect 58027 24160 58072 24188
rect 58066 24148 58072 24160
rect 58124 24148 58130 24200
rect 54812 24092 55720 24120
rect 54812 24080 54818 24092
rect 56870 24080 56876 24132
rect 56928 24120 56934 24132
rect 57977 24123 58035 24129
rect 57977 24120 57989 24123
rect 56928 24092 57989 24120
rect 56928 24080 56934 24092
rect 57977 24089 57989 24092
rect 58023 24089 58035 24123
rect 57977 24083 58035 24089
rect 27617 24055 27675 24061
rect 27617 24021 27629 24055
rect 27663 24052 27675 24055
rect 27798 24052 27804 24064
rect 27663 24024 27804 24052
rect 27663 24021 27675 24024
rect 27617 24015 27675 24021
rect 27798 24012 27804 24024
rect 27856 24012 27862 24064
rect 35621 24055 35679 24061
rect 35621 24021 35633 24055
rect 35667 24052 35679 24055
rect 39206 24052 39212 24064
rect 35667 24024 39212 24052
rect 35667 24021 35679 24024
rect 35621 24015 35679 24021
rect 39206 24012 39212 24024
rect 39264 24012 39270 24064
rect 40218 24012 40224 24064
rect 40276 24012 40282 24064
rect 44818 24012 44824 24064
rect 44876 24052 44882 24064
rect 45189 24055 45247 24061
rect 45189 24052 45201 24055
rect 44876 24024 45201 24052
rect 44876 24012 44882 24024
rect 45189 24021 45201 24024
rect 45235 24021 45247 24055
rect 46842 24052 46848 24064
rect 46803 24024 46848 24052
rect 45189 24015 45247 24021
rect 46842 24012 46848 24024
rect 46900 24012 46906 24064
rect 52825 24055 52883 24061
rect 52825 24021 52837 24055
rect 52871 24052 52883 24055
rect 56318 24052 56324 24064
rect 52871 24024 56324 24052
rect 52871 24021 52883 24024
rect 52825 24015 52883 24021
rect 56318 24012 56324 24024
rect 56376 24012 56382 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 28718 23808 28724 23860
rect 28776 23848 28782 23860
rect 28813 23851 28871 23857
rect 28813 23848 28825 23851
rect 28776 23820 28825 23848
rect 28776 23808 28782 23820
rect 28813 23817 28825 23820
rect 28859 23817 28871 23851
rect 31570 23848 31576 23860
rect 31531 23820 31576 23848
rect 28813 23811 28871 23817
rect 31570 23808 31576 23820
rect 31628 23808 31634 23860
rect 34977 23851 35035 23857
rect 34977 23817 34989 23851
rect 35023 23848 35035 23851
rect 35250 23848 35256 23860
rect 35023 23820 35256 23848
rect 35023 23817 35035 23820
rect 34977 23811 35035 23817
rect 35250 23808 35256 23820
rect 35308 23808 35314 23860
rect 36354 23848 36360 23860
rect 36315 23820 36360 23848
rect 36354 23808 36360 23820
rect 36412 23808 36418 23860
rect 38746 23848 38752 23860
rect 38707 23820 38752 23848
rect 38746 23808 38752 23820
rect 38804 23808 38810 23860
rect 39942 23848 39948 23860
rect 39903 23820 39948 23848
rect 39942 23808 39948 23820
rect 40000 23808 40006 23860
rect 40218 23808 40224 23860
rect 40276 23848 40282 23860
rect 42886 23848 42892 23860
rect 40276 23820 41000 23848
rect 40276 23808 40282 23820
rect 30558 23740 30564 23792
rect 30616 23780 30622 23792
rect 36446 23780 36452 23792
rect 30616 23752 31616 23780
rect 30616 23740 30622 23752
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23712 1918 23724
rect 2317 23715 2375 23721
rect 2317 23712 2329 23715
rect 1912 23684 2329 23712
rect 1912 23672 1918 23684
rect 2317 23681 2329 23684
rect 2363 23681 2375 23715
rect 2317 23675 2375 23681
rect 25038 23672 25044 23724
rect 25096 23672 25102 23724
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23712 25651 23715
rect 27522 23712 27528 23724
rect 25639 23684 27528 23712
rect 25639 23681 25651 23684
rect 25593 23675 25651 23681
rect 27522 23672 27528 23684
rect 27580 23672 27586 23724
rect 27798 23712 27804 23724
rect 27759 23684 27804 23712
rect 27798 23672 27804 23684
rect 27856 23672 27862 23724
rect 27982 23712 27988 23724
rect 27943 23684 27988 23712
rect 27982 23672 27988 23684
rect 28040 23672 28046 23724
rect 30190 23712 30196 23724
rect 30151 23684 30196 23712
rect 30190 23672 30196 23684
rect 30248 23672 30254 23724
rect 31588 23721 31616 23752
rect 35268 23752 36452 23780
rect 35268 23721 35296 23752
rect 36446 23740 36452 23752
rect 36504 23740 36510 23792
rect 38470 23740 38476 23792
rect 38528 23780 38534 23792
rect 38933 23783 38991 23789
rect 38933 23780 38945 23783
rect 38528 23752 38945 23780
rect 38528 23740 38534 23752
rect 38933 23749 38945 23752
rect 38979 23749 38991 23783
rect 38933 23743 38991 23749
rect 31389 23715 31447 23721
rect 31389 23681 31401 23715
rect 31435 23681 31447 23715
rect 31389 23675 31447 23681
rect 31573 23715 31631 23721
rect 31573 23681 31585 23715
rect 31619 23681 31631 23715
rect 31573 23675 31631 23681
rect 35253 23715 35311 23721
rect 35253 23681 35265 23715
rect 35299 23681 35311 23715
rect 35894 23712 35900 23724
rect 35855 23684 35900 23712
rect 35253 23675 35311 23681
rect 24394 23604 24400 23656
rect 24452 23644 24458 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 24452 23616 24593 23644
rect 24452 23604 24458 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 30009 23647 30067 23653
rect 30009 23613 30021 23647
rect 30055 23644 30067 23647
rect 31294 23644 31300 23656
rect 30055 23616 31300 23644
rect 30055 23613 30067 23616
rect 30009 23607 30067 23613
rect 31294 23604 31300 23616
rect 31352 23644 31358 23656
rect 31404 23644 31432 23675
rect 35894 23672 35900 23684
rect 35952 23712 35958 23724
rect 36357 23715 36415 23721
rect 36357 23712 36369 23715
rect 35952 23684 36369 23712
rect 35952 23672 35958 23684
rect 36357 23681 36369 23684
rect 36403 23681 36415 23715
rect 36357 23675 36415 23681
rect 36541 23715 36599 23721
rect 36541 23681 36553 23715
rect 36587 23681 36599 23715
rect 39114 23712 39120 23724
rect 39075 23684 39120 23712
rect 36541 23675 36599 23681
rect 31352 23616 31432 23644
rect 31352 23604 31358 23616
rect 34514 23604 34520 23656
rect 34572 23644 34578 23656
rect 34977 23647 35035 23653
rect 34977 23644 34989 23647
rect 34572 23616 34989 23644
rect 34572 23604 34578 23616
rect 34977 23613 34989 23616
rect 35023 23644 35035 23647
rect 36556 23644 36584 23675
rect 39114 23672 39120 23684
rect 39172 23672 39178 23724
rect 40218 23672 40224 23724
rect 40276 23712 40282 23724
rect 40405 23715 40463 23721
rect 40276 23684 40321 23712
rect 40276 23672 40282 23684
rect 40405 23681 40417 23715
rect 40451 23712 40463 23715
rect 40586 23712 40592 23724
rect 40451 23684 40592 23712
rect 40451 23681 40463 23684
rect 40405 23675 40463 23681
rect 40586 23672 40592 23684
rect 40644 23672 40650 23724
rect 40972 23721 41000 23820
rect 42628 23820 42892 23848
rect 40957 23715 41015 23721
rect 40957 23681 40969 23715
rect 41003 23681 41015 23715
rect 40957 23675 41015 23681
rect 41141 23715 41199 23721
rect 41141 23681 41153 23715
rect 41187 23712 41199 23715
rect 41230 23712 41236 23724
rect 41187 23684 41236 23712
rect 41187 23681 41199 23684
rect 41141 23675 41199 23681
rect 40126 23644 40132 23656
rect 35023 23616 36584 23644
rect 40087 23616 40132 23644
rect 35023 23613 35035 23616
rect 34977 23607 35035 23613
rect 40126 23604 40132 23616
rect 40184 23604 40190 23656
rect 40313 23647 40371 23653
rect 40313 23613 40325 23647
rect 40359 23644 40371 23647
rect 41156 23644 41184 23675
rect 41230 23672 41236 23684
rect 41288 23672 41294 23724
rect 42628 23721 42656 23820
rect 42886 23808 42892 23820
rect 42944 23848 42950 23860
rect 43898 23848 43904 23860
rect 42944 23820 43904 23848
rect 42944 23808 42950 23820
rect 43898 23808 43904 23820
rect 43956 23808 43962 23860
rect 44637 23851 44695 23857
rect 44637 23817 44649 23851
rect 44683 23848 44695 23851
rect 45925 23851 45983 23857
rect 44683 23820 45416 23848
rect 44683 23817 44695 23820
rect 44637 23811 44695 23817
rect 43438 23740 43444 23792
rect 43496 23780 43502 23792
rect 43496 23752 45232 23780
rect 43496 23740 43502 23752
rect 42613 23715 42671 23721
rect 42613 23681 42625 23715
rect 42659 23681 42671 23715
rect 42613 23675 42671 23681
rect 42797 23715 42855 23721
rect 42797 23681 42809 23715
rect 42843 23681 42855 23715
rect 42797 23675 42855 23681
rect 43901 23715 43959 23721
rect 43901 23681 43913 23715
rect 43947 23712 43959 23715
rect 44174 23712 44180 23724
rect 43947 23684 44180 23712
rect 43947 23681 43959 23684
rect 43901 23675 43959 23681
rect 40359 23616 41184 23644
rect 42812 23644 42840 23675
rect 44174 23672 44180 23684
rect 44232 23672 44238 23724
rect 44450 23712 44456 23724
rect 44411 23684 44456 23712
rect 44450 23672 44456 23684
rect 44508 23672 44514 23724
rect 45204 23721 45232 23752
rect 45388 23721 45416 23820
rect 45925 23817 45937 23851
rect 45971 23848 45983 23851
rect 46014 23848 46020 23860
rect 45971 23820 46020 23848
rect 45971 23817 45983 23820
rect 45925 23811 45983 23817
rect 46014 23808 46020 23820
rect 46072 23808 46078 23860
rect 46842 23808 46848 23860
rect 46900 23848 46906 23860
rect 47965 23851 48023 23857
rect 47965 23848 47977 23851
rect 46900 23820 47977 23848
rect 46900 23808 46906 23820
rect 47965 23817 47977 23820
rect 48011 23817 48023 23851
rect 47965 23811 48023 23817
rect 48133 23851 48191 23857
rect 48133 23817 48145 23851
rect 48179 23848 48191 23851
rect 49878 23848 49884 23860
rect 48179 23820 49740 23848
rect 49839 23820 49884 23848
rect 48179 23817 48191 23820
rect 48133 23811 48191 23817
rect 46198 23740 46204 23792
rect 46256 23780 46262 23792
rect 47765 23783 47823 23789
rect 47765 23780 47777 23783
rect 46256 23752 47777 23780
rect 46256 23740 46262 23752
rect 47765 23749 47777 23752
rect 47811 23749 47823 23783
rect 48590 23780 48596 23792
rect 48551 23752 48596 23780
rect 47765 23743 47823 23749
rect 48590 23740 48596 23752
rect 48648 23740 48654 23792
rect 48809 23783 48867 23789
rect 48809 23749 48821 23783
rect 48855 23780 48867 23783
rect 48958 23780 48964 23792
rect 48855 23752 48964 23780
rect 48855 23749 48867 23752
rect 48809 23743 48867 23749
rect 48958 23740 48964 23752
rect 49016 23740 49022 23792
rect 49712 23724 49740 23820
rect 49878 23808 49884 23820
rect 49936 23808 49942 23860
rect 50798 23848 50804 23860
rect 50759 23820 50804 23848
rect 50798 23808 50804 23820
rect 50856 23808 50862 23860
rect 53098 23848 53104 23860
rect 53059 23820 53104 23848
rect 53098 23808 53104 23820
rect 53156 23808 53162 23860
rect 54202 23848 54208 23860
rect 54163 23820 54208 23848
rect 54202 23808 54208 23820
rect 54260 23808 54266 23860
rect 56410 23848 56416 23860
rect 56371 23820 56416 23848
rect 56410 23808 56416 23820
rect 56468 23808 56474 23860
rect 58158 23848 58164 23860
rect 58119 23820 58164 23848
rect 58158 23808 58164 23820
rect 58216 23808 58222 23860
rect 50062 23740 50068 23792
rect 50120 23780 50126 23792
rect 50433 23783 50491 23789
rect 50433 23780 50445 23783
rect 50120 23752 50445 23780
rect 50120 23740 50126 23752
rect 50433 23749 50445 23752
rect 50479 23780 50491 23783
rect 50479 23752 51304 23780
rect 50479 23749 50491 23752
rect 50433 23743 50491 23749
rect 45189 23715 45247 23721
rect 45189 23681 45201 23715
rect 45235 23681 45247 23715
rect 45189 23675 45247 23681
rect 45373 23715 45431 23721
rect 45373 23681 45385 23715
rect 45419 23681 45431 23715
rect 46658 23712 46664 23724
rect 46619 23684 46664 23712
rect 45373 23675 45431 23681
rect 45281 23647 45339 23653
rect 45281 23644 45293 23647
rect 42812 23616 45293 23644
rect 40359 23613 40371 23616
rect 40313 23607 40371 23613
rect 45281 23613 45293 23616
rect 45327 23613 45339 23647
rect 45388 23644 45416 23675
rect 46658 23672 46664 23684
rect 46716 23672 46722 23724
rect 46750 23672 46756 23724
rect 46808 23712 46814 23724
rect 46934 23712 46940 23724
rect 46808 23684 46853 23712
rect 46895 23684 46940 23712
rect 46808 23672 46814 23684
rect 46934 23672 46940 23684
rect 46992 23712 46998 23724
rect 47302 23712 47308 23724
rect 46992 23684 47308 23712
rect 46992 23672 46998 23684
rect 47302 23672 47308 23684
rect 47360 23672 47366 23724
rect 49694 23712 49700 23724
rect 49607 23684 49700 23712
rect 49694 23672 49700 23684
rect 49752 23672 49758 23724
rect 49970 23672 49976 23724
rect 50028 23712 50034 23724
rect 51276 23721 51304 23752
rect 51994 23740 52000 23792
rect 52052 23780 52058 23792
rect 52365 23783 52423 23789
rect 52365 23780 52377 23783
rect 52052 23752 52377 23780
rect 52052 23740 52058 23752
rect 52365 23749 52377 23752
rect 52411 23749 52423 23783
rect 52365 23743 52423 23749
rect 50617 23715 50675 23721
rect 50617 23712 50629 23715
rect 50028 23684 50629 23712
rect 50028 23672 50034 23684
rect 50617 23681 50629 23684
rect 50663 23681 50675 23715
rect 50617 23675 50675 23681
rect 51261 23715 51319 23721
rect 51261 23681 51273 23715
rect 51307 23681 51319 23715
rect 51261 23675 51319 23681
rect 51445 23715 51503 23721
rect 51445 23681 51457 23715
rect 51491 23712 51503 23715
rect 51626 23712 51632 23724
rect 51491 23684 51632 23712
rect 51491 23681 51503 23684
rect 51445 23675 51503 23681
rect 51626 23672 51632 23684
rect 51684 23672 51690 23724
rect 52086 23712 52092 23724
rect 52047 23684 52092 23712
rect 52086 23672 52092 23684
rect 52144 23672 52150 23724
rect 52178 23672 52184 23724
rect 52236 23712 52242 23724
rect 53006 23712 53012 23724
rect 52236 23684 52281 23712
rect 52967 23684 53012 23712
rect 52236 23672 52242 23684
rect 53006 23672 53012 23684
rect 53064 23672 53070 23724
rect 53193 23715 53251 23721
rect 53193 23681 53205 23715
rect 53239 23712 53251 23715
rect 53282 23712 53288 23724
rect 53239 23684 53288 23712
rect 53239 23681 53251 23684
rect 53193 23675 53251 23681
rect 53282 23672 53288 23684
rect 53340 23672 53346 23724
rect 53834 23712 53840 23724
rect 53795 23684 53840 23712
rect 53834 23672 53840 23684
rect 53892 23672 53898 23724
rect 56318 23712 56324 23724
rect 56279 23684 56324 23712
rect 56318 23672 56324 23684
rect 56376 23672 56382 23724
rect 56410 23672 56416 23724
rect 56468 23712 56474 23724
rect 56505 23715 56563 23721
rect 56505 23712 56517 23715
rect 56468 23684 56517 23712
rect 56468 23672 56474 23684
rect 56505 23681 56517 23684
rect 56551 23681 56563 23715
rect 58158 23712 58164 23724
rect 56505 23675 56563 23681
rect 56980 23684 58164 23712
rect 48590 23644 48596 23656
rect 45388 23616 48596 23644
rect 45281 23607 45339 23613
rect 48590 23604 48596 23616
rect 48648 23604 48654 23656
rect 49418 23644 49424 23656
rect 49379 23616 49424 23644
rect 49418 23604 49424 23616
rect 49476 23604 49482 23656
rect 53926 23644 53932 23656
rect 53887 23616 53932 23644
rect 53926 23604 53932 23616
rect 53984 23604 53990 23656
rect 56980 23644 57008 23684
rect 58158 23672 58164 23684
rect 58216 23712 58222 23724
rect 58345 23715 58403 23721
rect 58345 23712 58357 23715
rect 58216 23684 58357 23712
rect 58216 23672 58222 23684
rect 58345 23681 58357 23684
rect 58391 23681 58403 23715
rect 58345 23675 58403 23681
rect 55186 23616 57008 23644
rect 57057 23647 57115 23653
rect 30377 23579 30435 23585
rect 30377 23545 30389 23579
rect 30423 23576 30435 23579
rect 55186 23576 55214 23616
rect 57057 23613 57069 23647
rect 57103 23644 57115 23647
rect 57422 23644 57428 23656
rect 57103 23616 57428 23644
rect 57103 23613 57115 23616
rect 57057 23607 57115 23613
rect 57422 23604 57428 23616
rect 57480 23604 57486 23656
rect 30423 23548 55214 23576
rect 30423 23545 30435 23548
rect 30377 23539 30435 23545
rect 56870 23536 56876 23588
rect 56928 23576 56934 23588
rect 57333 23579 57391 23585
rect 57333 23576 57345 23579
rect 56928 23548 57345 23576
rect 56928 23536 56934 23548
rect 57333 23545 57345 23548
rect 57379 23545 57391 23579
rect 57333 23539 57391 23545
rect 1670 23508 1676 23520
rect 1631 23480 1676 23508
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 35161 23511 35219 23517
rect 35161 23477 35173 23511
rect 35207 23508 35219 23511
rect 35805 23511 35863 23517
rect 35805 23508 35817 23511
rect 35207 23480 35817 23508
rect 35207 23477 35219 23480
rect 35161 23471 35219 23477
rect 35805 23477 35817 23480
rect 35851 23477 35863 23511
rect 35805 23471 35863 23477
rect 40862 23468 40868 23520
rect 40920 23508 40926 23520
rect 41049 23511 41107 23517
rect 41049 23508 41061 23511
rect 40920 23480 41061 23508
rect 40920 23468 40926 23480
rect 41049 23477 41061 23480
rect 41095 23477 41107 23511
rect 41690 23508 41696 23520
rect 41651 23480 41696 23508
rect 41049 23471 41107 23477
rect 41690 23468 41696 23480
rect 41748 23468 41754 23520
rect 41966 23468 41972 23520
rect 42024 23508 42030 23520
rect 42705 23511 42763 23517
rect 42705 23508 42717 23511
rect 42024 23480 42717 23508
rect 42024 23468 42030 23480
rect 42705 23477 42717 23480
rect 42751 23477 42763 23511
rect 42705 23471 42763 23477
rect 43809 23511 43867 23517
rect 43809 23477 43821 23511
rect 43855 23508 43867 23511
rect 44450 23508 44456 23520
rect 43855 23480 44456 23508
rect 43855 23477 43867 23480
rect 43809 23471 43867 23477
rect 44450 23468 44456 23480
rect 44508 23468 44514 23520
rect 47121 23511 47179 23517
rect 47121 23477 47133 23511
rect 47167 23508 47179 23511
rect 47949 23511 48007 23517
rect 47949 23508 47961 23511
rect 47167 23480 47961 23508
rect 47167 23477 47179 23480
rect 47121 23471 47179 23477
rect 47949 23477 47961 23480
rect 47995 23477 48007 23511
rect 47949 23471 48007 23477
rect 48682 23468 48688 23520
rect 48740 23508 48746 23520
rect 48777 23511 48835 23517
rect 48777 23508 48789 23511
rect 48740 23480 48789 23508
rect 48740 23468 48746 23480
rect 48777 23477 48789 23480
rect 48823 23477 48835 23511
rect 48777 23471 48835 23477
rect 48961 23511 49019 23517
rect 48961 23477 48973 23511
rect 49007 23508 49019 23511
rect 49234 23508 49240 23520
rect 49007 23480 49240 23508
rect 49007 23477 49019 23480
rect 48961 23471 49019 23477
rect 49234 23468 49240 23480
rect 49292 23468 49298 23520
rect 49513 23511 49571 23517
rect 49513 23477 49525 23511
rect 49559 23508 49571 23511
rect 49786 23508 49792 23520
rect 49559 23480 49792 23508
rect 49559 23477 49571 23480
rect 49513 23471 49571 23477
rect 49786 23468 49792 23480
rect 49844 23468 49850 23520
rect 51629 23511 51687 23517
rect 51629 23477 51641 23511
rect 51675 23508 51687 23511
rect 51902 23508 51908 23520
rect 51675 23480 51908 23508
rect 51675 23477 51687 23480
rect 51629 23471 51687 23477
rect 51902 23468 51908 23480
rect 51960 23468 51966 23520
rect 52365 23511 52423 23517
rect 52365 23477 52377 23511
rect 52411 23508 52423 23511
rect 52454 23508 52460 23520
rect 52411 23480 52460 23508
rect 52411 23477 52423 23480
rect 52365 23471 52423 23477
rect 52454 23468 52460 23480
rect 52512 23468 52518 23520
rect 57517 23511 57575 23517
rect 57517 23477 57529 23511
rect 57563 23508 57575 23511
rect 57790 23508 57796 23520
rect 57563 23480 57796 23508
rect 57563 23477 57575 23480
rect 57517 23471 57575 23477
rect 57790 23468 57796 23480
rect 57848 23468 57854 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 27522 23264 27528 23316
rect 27580 23304 27586 23316
rect 28445 23307 28503 23313
rect 28445 23304 28457 23307
rect 27580 23276 28457 23304
rect 27580 23264 27586 23276
rect 28445 23273 28457 23276
rect 28491 23273 28503 23307
rect 28445 23267 28503 23273
rect 29733 23307 29791 23313
rect 29733 23273 29745 23307
rect 29779 23304 29791 23307
rect 30190 23304 30196 23316
rect 29779 23276 30196 23304
rect 29779 23273 29791 23276
rect 29733 23267 29791 23273
rect 30190 23264 30196 23276
rect 30248 23264 30254 23316
rect 34241 23307 34299 23313
rect 34241 23273 34253 23307
rect 34287 23304 34299 23307
rect 34514 23304 34520 23316
rect 34287 23276 34520 23304
rect 34287 23273 34299 23276
rect 34241 23267 34299 23273
rect 34514 23264 34520 23276
rect 34572 23264 34578 23316
rect 35345 23307 35403 23313
rect 35345 23273 35357 23307
rect 35391 23304 35403 23307
rect 35894 23304 35900 23316
rect 35391 23276 35900 23304
rect 35391 23273 35403 23276
rect 35345 23267 35403 23273
rect 35894 23264 35900 23276
rect 35952 23264 35958 23316
rect 38470 23264 38476 23316
rect 38528 23304 38534 23316
rect 38565 23307 38623 23313
rect 38565 23304 38577 23307
rect 38528 23276 38577 23304
rect 38528 23264 38534 23276
rect 38565 23273 38577 23276
rect 38611 23273 38623 23307
rect 38565 23267 38623 23273
rect 39025 23307 39083 23313
rect 39025 23273 39037 23307
rect 39071 23304 39083 23307
rect 39114 23304 39120 23316
rect 39071 23276 39120 23304
rect 39071 23273 39083 23276
rect 39025 23267 39083 23273
rect 39114 23264 39120 23276
rect 39172 23264 39178 23316
rect 43438 23304 43444 23316
rect 43399 23276 43444 23304
rect 43438 23264 43444 23276
rect 43496 23264 43502 23316
rect 45649 23307 45707 23313
rect 45649 23273 45661 23307
rect 45695 23304 45707 23307
rect 45738 23304 45744 23316
rect 45695 23276 45744 23304
rect 45695 23273 45707 23276
rect 45649 23267 45707 23273
rect 45738 23264 45744 23276
rect 45796 23264 45802 23316
rect 46477 23307 46535 23313
rect 46477 23273 46489 23307
rect 46523 23304 46535 23307
rect 46658 23304 46664 23316
rect 46523 23276 46664 23304
rect 46523 23273 46535 23276
rect 46477 23267 46535 23273
rect 46658 23264 46664 23276
rect 46716 23264 46722 23316
rect 48961 23307 49019 23313
rect 48961 23273 48973 23307
rect 49007 23304 49019 23307
rect 49142 23304 49148 23316
rect 49007 23276 49148 23304
rect 49007 23273 49019 23276
rect 48961 23267 49019 23273
rect 49142 23264 49148 23276
rect 49200 23264 49206 23316
rect 49789 23307 49847 23313
rect 49789 23273 49801 23307
rect 49835 23304 49847 23307
rect 50154 23304 50160 23316
rect 49835 23276 50160 23304
rect 49835 23273 49847 23276
rect 49789 23267 49847 23273
rect 50154 23264 50160 23276
rect 50212 23264 50218 23316
rect 52086 23304 52092 23316
rect 52047 23276 52092 23304
rect 52086 23264 52092 23276
rect 52144 23264 52150 23316
rect 52273 23307 52331 23313
rect 52273 23273 52285 23307
rect 52319 23304 52331 23307
rect 53190 23304 53196 23316
rect 52319 23276 53196 23304
rect 52319 23273 52331 23276
rect 52273 23267 52331 23273
rect 53190 23264 53196 23276
rect 53248 23264 53254 23316
rect 53282 23264 53288 23316
rect 53340 23304 53346 23316
rect 53561 23307 53619 23313
rect 53561 23304 53573 23307
rect 53340 23276 53573 23304
rect 53340 23264 53346 23276
rect 53561 23273 53573 23276
rect 53607 23273 53619 23307
rect 53561 23267 53619 23273
rect 53745 23307 53803 23313
rect 53745 23273 53757 23307
rect 53791 23304 53803 23307
rect 53834 23304 53840 23316
rect 53791 23276 53840 23304
rect 53791 23273 53803 23276
rect 53745 23267 53803 23273
rect 53834 23264 53840 23276
rect 53892 23264 53898 23316
rect 57606 23304 57612 23316
rect 57567 23276 57612 23304
rect 57606 23264 57612 23276
rect 57664 23264 57670 23316
rect 58066 23264 58072 23316
rect 58124 23304 58130 23316
rect 58253 23307 58311 23313
rect 58253 23304 58265 23307
rect 58124 23276 58265 23304
rect 58124 23264 58130 23276
rect 58253 23273 58265 23276
rect 58299 23273 58311 23307
rect 58253 23267 58311 23273
rect 28626 23236 28632 23248
rect 28539 23208 28632 23236
rect 28626 23196 28632 23208
rect 28684 23236 28690 23248
rect 31018 23236 31024 23248
rect 28684 23208 31024 23236
rect 28684 23196 28690 23208
rect 31018 23196 31024 23208
rect 31076 23196 31082 23248
rect 44637 23239 44695 23245
rect 35360 23208 37412 23236
rect 26145 23171 26203 23177
rect 26145 23168 26157 23171
rect 23584 23140 26157 23168
rect 22830 23060 22836 23112
rect 22888 23100 22894 23112
rect 23109 23103 23167 23109
rect 23109 23100 23121 23103
rect 22888 23072 23121 23100
rect 22888 23060 22894 23072
rect 23109 23069 23121 23072
rect 23155 23069 23167 23103
rect 23109 23063 23167 23069
rect 23382 23060 23388 23112
rect 23440 23100 23446 23112
rect 23584 23109 23612 23140
rect 26145 23137 26157 23140
rect 26191 23137 26203 23171
rect 26145 23131 26203 23137
rect 31113 23171 31171 23177
rect 31113 23137 31125 23171
rect 31159 23168 31171 23171
rect 32490 23168 32496 23180
rect 31159 23140 32496 23168
rect 31159 23137 31171 23140
rect 31113 23131 31171 23137
rect 32490 23128 32496 23140
rect 32548 23128 32554 23180
rect 35360 23112 35388 23208
rect 36357 23171 36415 23177
rect 36357 23137 36369 23171
rect 36403 23168 36415 23171
rect 36446 23168 36452 23180
rect 36403 23140 36452 23168
rect 36403 23137 36415 23140
rect 36357 23131 36415 23137
rect 36446 23128 36452 23140
rect 36504 23128 36510 23180
rect 37384 23177 37412 23208
rect 44637 23205 44649 23239
rect 44683 23236 44695 23239
rect 45002 23236 45008 23248
rect 44683 23208 45008 23236
rect 44683 23205 44695 23208
rect 44637 23199 44695 23205
rect 45002 23196 45008 23208
rect 45060 23196 45066 23248
rect 45281 23239 45339 23245
rect 45281 23205 45293 23239
rect 45327 23236 45339 23239
rect 45554 23236 45560 23248
rect 45327 23208 45560 23236
rect 45327 23205 45339 23208
rect 45281 23199 45339 23205
rect 45554 23196 45560 23208
rect 45612 23196 45618 23248
rect 49694 23236 49700 23248
rect 49655 23208 49700 23236
rect 49694 23196 49700 23208
rect 49752 23196 49758 23248
rect 49970 23196 49976 23248
rect 50028 23236 50034 23248
rect 50341 23239 50399 23245
rect 50341 23236 50353 23239
rect 50028 23208 50353 23236
rect 50028 23196 50034 23208
rect 50341 23205 50353 23208
rect 50387 23205 50399 23239
rect 50341 23199 50399 23205
rect 56045 23239 56103 23245
rect 56045 23205 56057 23239
rect 56091 23236 56103 23239
rect 56134 23236 56140 23248
rect 56091 23208 56140 23236
rect 56091 23205 56103 23208
rect 56045 23199 56103 23205
rect 56134 23196 56140 23208
rect 56192 23196 56198 23248
rect 36633 23171 36691 23177
rect 36633 23137 36645 23171
rect 36679 23137 36691 23171
rect 36633 23131 36691 23137
rect 37369 23171 37427 23177
rect 37369 23137 37381 23171
rect 37415 23168 37427 23171
rect 37458 23168 37464 23180
rect 37415 23140 37464 23168
rect 37415 23137 37427 23140
rect 37369 23131 37427 23137
rect 23569 23103 23627 23109
rect 23569 23100 23581 23103
rect 23440 23072 23581 23100
rect 23440 23060 23446 23072
rect 23569 23069 23581 23072
rect 23615 23069 23627 23103
rect 23569 23063 23627 23069
rect 26053 23103 26111 23109
rect 26053 23069 26065 23103
rect 26099 23100 26111 23103
rect 26234 23100 26240 23112
rect 26099 23072 26240 23100
rect 26099 23069 26111 23072
rect 26053 23063 26111 23069
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 26694 23100 26700 23112
rect 26655 23072 26700 23100
rect 26694 23060 26700 23072
rect 26752 23060 26758 23112
rect 27062 23100 27068 23112
rect 27023 23072 27068 23100
rect 27062 23060 27068 23072
rect 27120 23060 27126 23112
rect 27433 23103 27491 23109
rect 27433 23069 27445 23103
rect 27479 23100 27491 23103
rect 27522 23100 27528 23112
rect 27479 23072 27528 23100
rect 27479 23069 27491 23072
rect 27433 23063 27491 23069
rect 27522 23060 27528 23072
rect 27580 23060 27586 23112
rect 27982 23100 27988 23112
rect 27943 23072 27988 23100
rect 27982 23060 27988 23072
rect 28040 23060 28046 23112
rect 28994 23060 29000 23112
rect 29052 23100 29058 23112
rect 29917 23103 29975 23109
rect 29917 23100 29929 23103
rect 29052 23072 29929 23100
rect 29052 23060 29058 23072
rect 29917 23069 29929 23072
rect 29963 23069 29975 23103
rect 29917 23063 29975 23069
rect 30193 23103 30251 23109
rect 30193 23069 30205 23103
rect 30239 23100 30251 23103
rect 30558 23100 30564 23112
rect 30239 23072 30564 23100
rect 30239 23069 30251 23072
rect 30193 23063 30251 23069
rect 30558 23060 30564 23072
rect 30616 23060 30622 23112
rect 30742 23100 30748 23112
rect 30703 23072 30748 23100
rect 30742 23060 30748 23072
rect 30800 23060 30806 23112
rect 31021 23103 31079 23109
rect 31021 23069 31033 23103
rect 31067 23100 31079 23103
rect 31662 23100 31668 23112
rect 31067 23072 31668 23100
rect 31067 23069 31079 23072
rect 31021 23063 31079 23069
rect 31662 23060 31668 23072
rect 31720 23060 31726 23112
rect 31757 23103 31815 23109
rect 31757 23069 31769 23103
rect 31803 23069 31815 23103
rect 31757 23063 31815 23069
rect 31849 23103 31907 23109
rect 31849 23069 31861 23103
rect 31895 23069 31907 23103
rect 31849 23063 31907 23069
rect 31941 23103 31999 23109
rect 31941 23069 31953 23103
rect 31987 23100 31999 23103
rect 32122 23100 32128 23112
rect 31987 23072 32128 23100
rect 31987 23069 31999 23072
rect 31941 23063 31999 23069
rect 28534 22992 28540 23044
rect 28592 23032 28598 23044
rect 28905 23035 28963 23041
rect 28905 23032 28917 23035
rect 28592 23004 28917 23032
rect 28592 22992 28598 23004
rect 28905 23001 28917 23004
rect 28951 23032 28963 23035
rect 29454 23032 29460 23044
rect 28951 23004 29460 23032
rect 28951 23001 28963 23004
rect 28905 22995 28963 23001
rect 29454 22992 29460 23004
rect 29512 22992 29518 23044
rect 30576 23032 30604 23060
rect 31772 23032 31800 23063
rect 30576 23004 31800 23032
rect 31864 22976 31892 23063
rect 32122 23060 32128 23072
rect 32180 23060 32186 23112
rect 34149 23103 34207 23109
rect 34149 23069 34161 23103
rect 34195 23069 34207 23103
rect 34149 23063 34207 23069
rect 34333 23103 34391 23109
rect 34333 23069 34345 23103
rect 34379 23100 34391 23103
rect 35161 23103 35219 23109
rect 35161 23100 35173 23103
rect 34379 23072 35173 23100
rect 34379 23069 34391 23072
rect 34333 23063 34391 23069
rect 35161 23069 35173 23072
rect 35207 23100 35219 23103
rect 35342 23100 35348 23112
rect 35207 23072 35348 23100
rect 35207 23069 35219 23072
rect 35161 23063 35219 23069
rect 34164 23032 34192 23063
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 36262 23100 36268 23112
rect 36223 23072 36268 23100
rect 36262 23060 36268 23072
rect 36320 23060 36326 23112
rect 36648 23100 36676 23131
rect 37458 23128 37464 23140
rect 37516 23128 37522 23180
rect 37645 23171 37703 23177
rect 37645 23137 37657 23171
rect 37691 23168 37703 23171
rect 41966 23168 41972 23180
rect 37691 23140 38424 23168
rect 41927 23140 41972 23168
rect 37691 23137 37703 23140
rect 37645 23131 37703 23137
rect 37274 23100 37280 23112
rect 36648 23072 37280 23100
rect 37274 23060 37280 23072
rect 37332 23060 37338 23112
rect 38102 23100 38108 23112
rect 38063 23072 38108 23100
rect 38102 23060 38108 23072
rect 38160 23060 38166 23112
rect 38197 23103 38255 23109
rect 38197 23069 38209 23103
rect 38243 23100 38255 23103
rect 38286 23100 38292 23112
rect 38243 23072 38292 23100
rect 38243 23069 38255 23072
rect 38197 23063 38255 23069
rect 38286 23060 38292 23072
rect 38344 23060 38350 23112
rect 38396 23109 38424 23140
rect 41966 23128 41972 23140
rect 42024 23128 42030 23180
rect 44358 23168 44364 23180
rect 44319 23140 44364 23168
rect 44358 23128 44364 23140
rect 44416 23128 44422 23180
rect 47673 23171 47731 23177
rect 47673 23168 47685 23171
rect 45572 23140 46336 23168
rect 45572 23112 45600 23140
rect 38381 23103 38439 23109
rect 38381 23069 38393 23103
rect 38427 23100 38439 23103
rect 39025 23103 39083 23109
rect 39025 23100 39037 23103
rect 38427 23072 39037 23100
rect 38427 23069 38439 23072
rect 38381 23063 38439 23069
rect 39025 23069 39037 23072
rect 39071 23069 39083 23103
rect 39025 23063 39083 23069
rect 39117 23103 39175 23109
rect 39117 23069 39129 23103
rect 39163 23069 39175 23103
rect 40494 23100 40500 23112
rect 40455 23072 40500 23100
rect 39117 23063 39175 23069
rect 34698 23032 34704 23044
rect 34164 23004 34704 23032
rect 34698 22992 34704 23004
rect 34756 23032 34762 23044
rect 34977 23035 35035 23041
rect 34977 23032 34989 23035
rect 34756 23004 34989 23032
rect 34756 22992 34762 23004
rect 34977 23001 34989 23004
rect 35023 23001 35035 23035
rect 36280 23032 36308 23060
rect 36722 23032 36728 23044
rect 36280 23004 36728 23032
rect 34977 22995 35035 23001
rect 36722 22992 36728 23004
rect 36780 22992 36786 23044
rect 38304 23032 38332 23060
rect 39132 23032 39160 23063
rect 40494 23060 40500 23072
rect 40552 23060 40558 23112
rect 40862 23100 40868 23112
rect 40823 23072 40868 23100
rect 40862 23060 40868 23072
rect 40920 23060 40926 23112
rect 41598 23060 41604 23112
rect 41656 23100 41662 23112
rect 41693 23103 41751 23109
rect 41693 23100 41705 23103
rect 41656 23072 41705 23100
rect 41656 23060 41662 23072
rect 41693 23069 41705 23072
rect 41739 23069 41751 23103
rect 44266 23100 44272 23112
rect 44227 23072 44272 23100
rect 41693 23063 41751 23069
rect 44266 23060 44272 23072
rect 44324 23060 44330 23112
rect 44634 23060 44640 23112
rect 44692 23060 44698 23112
rect 45554 23100 45560 23112
rect 45515 23072 45560 23100
rect 45554 23060 45560 23072
rect 45612 23060 45618 23112
rect 45649 23103 45707 23109
rect 45649 23069 45661 23103
rect 45695 23100 45707 23103
rect 46014 23100 46020 23112
rect 45695 23072 46020 23100
rect 45695 23069 45707 23072
rect 45649 23063 45707 23069
rect 46014 23060 46020 23072
rect 46072 23060 46078 23112
rect 46308 23109 46336 23140
rect 46676 23140 47685 23168
rect 46293 23103 46351 23109
rect 46293 23069 46305 23103
rect 46339 23069 46351 23103
rect 46293 23063 46351 23069
rect 38304 23004 39160 23032
rect 39301 23035 39359 23041
rect 39301 23001 39313 23035
rect 39347 23001 39359 23035
rect 39301 22995 39359 23001
rect 15930 22924 15936 22976
rect 15988 22964 15994 22976
rect 22741 22967 22799 22973
rect 22741 22964 22753 22967
rect 15988 22936 22753 22964
rect 15988 22924 15994 22936
rect 22741 22933 22753 22936
rect 22787 22933 22799 22967
rect 22741 22927 22799 22933
rect 30101 22967 30159 22973
rect 30101 22933 30113 22967
rect 30147 22964 30159 22967
rect 30282 22964 30288 22976
rect 30147 22936 30288 22964
rect 30147 22933 30159 22936
rect 30101 22927 30159 22933
rect 30282 22924 30288 22936
rect 30340 22924 30346 22976
rect 31846 22924 31852 22976
rect 31904 22924 31910 22976
rect 32125 22967 32183 22973
rect 32125 22933 32137 22967
rect 32171 22964 32183 22967
rect 33962 22964 33968 22976
rect 32171 22936 33968 22964
rect 32171 22933 32183 22936
rect 32125 22927 32183 22933
rect 33962 22924 33968 22936
rect 34020 22924 34026 22976
rect 38102 22924 38108 22976
rect 38160 22964 38166 22976
rect 39316 22964 39344 22995
rect 42426 22992 42432 23044
rect 42484 22992 42490 23044
rect 44652 23032 44680 23060
rect 46109 23035 46167 23041
rect 46109 23032 46121 23035
rect 44652 23004 46121 23032
rect 46109 23001 46121 23004
rect 46155 23032 46167 23035
rect 46676 23032 46704 23140
rect 47673 23137 47685 23140
rect 47719 23168 47731 23171
rect 48038 23168 48044 23180
rect 47719 23140 48044 23168
rect 47719 23137 47731 23140
rect 47673 23131 47731 23137
rect 48038 23128 48044 23140
rect 48096 23128 48102 23180
rect 48133 23171 48191 23177
rect 48133 23137 48145 23171
rect 48179 23137 48191 23171
rect 55582 23168 55588 23180
rect 55543 23140 55588 23168
rect 48133 23131 48191 23137
rect 46750 23060 46756 23112
rect 46808 23100 46814 23112
rect 47765 23103 47823 23109
rect 47765 23100 47777 23103
rect 46808 23072 47777 23100
rect 46808 23060 46814 23072
rect 47765 23069 47777 23072
rect 47811 23069 47823 23103
rect 48148 23100 48176 23131
rect 55582 23128 55588 23140
rect 55640 23128 55646 23180
rect 48682 23100 48688 23112
rect 48148 23072 48688 23100
rect 47765 23063 47823 23069
rect 48682 23060 48688 23072
rect 48740 23060 48746 23112
rect 48958 23100 48964 23112
rect 48919 23072 48964 23100
rect 48958 23060 48964 23072
rect 49016 23060 49022 23112
rect 49786 23060 49792 23112
rect 49844 23100 49850 23112
rect 52178 23100 52184 23112
rect 49844 23072 49889 23100
rect 51920 23072 52184 23100
rect 49844 23060 49850 23072
rect 46155 23004 46704 23032
rect 46155 23001 46167 23004
rect 46109 22995 46167 23001
rect 49418 22992 49424 23044
rect 49476 23032 49482 23044
rect 51920 23041 51948 23072
rect 52178 23060 52184 23072
rect 52236 23060 52242 23112
rect 55674 23100 55680 23112
rect 55635 23072 55680 23100
rect 55674 23060 55680 23072
rect 55732 23060 55738 23112
rect 58069 23103 58127 23109
rect 58069 23069 58081 23103
rect 58115 23069 58127 23103
rect 58250 23100 58256 23112
rect 58211 23072 58256 23100
rect 58069 23063 58127 23069
rect 49513 23035 49571 23041
rect 49513 23032 49525 23035
rect 49476 23004 49525 23032
rect 49476 22992 49482 23004
rect 49513 23001 49525 23004
rect 49559 23001 49571 23035
rect 51905 23035 51963 23041
rect 51905 23032 51917 23035
rect 49513 22995 49571 23001
rect 49620 23004 51917 23032
rect 38160 22936 39344 22964
rect 41233 22967 41291 22973
rect 38160 22924 38166 22936
rect 41233 22933 41245 22967
rect 41279 22964 41291 22967
rect 44542 22964 44548 22976
rect 41279 22936 44548 22964
rect 41279 22933 41291 22936
rect 41233 22927 41291 22933
rect 44542 22924 44548 22936
rect 44600 22924 44606 22976
rect 48590 22924 48596 22976
rect 48648 22964 48654 22976
rect 48777 22967 48835 22973
rect 48777 22964 48789 22967
rect 48648 22936 48789 22964
rect 48648 22924 48654 22936
rect 48777 22933 48789 22936
rect 48823 22964 48835 22967
rect 49620 22964 49648 23004
rect 51905 23001 51917 23004
rect 51951 23001 51963 23035
rect 51905 22995 51963 23001
rect 53006 22992 53012 23044
rect 53064 23032 53070 23044
rect 53190 23032 53196 23044
rect 53064 23004 53196 23032
rect 53064 22992 53070 23004
rect 53190 22992 53196 23004
rect 53248 23032 53254 23044
rect 53377 23035 53435 23041
rect 53377 23032 53389 23035
rect 53248 23004 53389 23032
rect 53248 22992 53254 23004
rect 53377 23001 53389 23004
rect 53423 23001 53435 23035
rect 53377 22995 53435 23001
rect 53593 23035 53651 23041
rect 53593 23001 53605 23035
rect 53639 23032 53651 23035
rect 54662 23032 54668 23044
rect 53639 23004 54668 23032
rect 53639 23001 53651 23004
rect 53593 22995 53651 23001
rect 54662 22992 54668 23004
rect 54720 22992 54726 23044
rect 56962 22992 56968 23044
rect 57020 23032 57026 23044
rect 57241 23035 57299 23041
rect 57241 23032 57253 23035
rect 57020 23004 57253 23032
rect 57020 22992 57026 23004
rect 57241 23001 57253 23004
rect 57287 23001 57299 23035
rect 57422 23032 57428 23044
rect 57383 23004 57428 23032
rect 57241 22995 57299 23001
rect 57422 22992 57428 23004
rect 57480 23032 57486 23044
rect 58084 23032 58112 23063
rect 58250 23060 58256 23072
rect 58308 23060 58314 23112
rect 57480 23004 58112 23032
rect 57480 22992 57486 23004
rect 48823 22936 49648 22964
rect 48823 22933 48835 22936
rect 48777 22927 48835 22933
rect 51994 22924 52000 22976
rect 52052 22964 52058 22976
rect 52105 22967 52163 22973
rect 52105 22964 52117 22967
rect 52052 22936 52117 22964
rect 52052 22924 52058 22936
rect 52105 22933 52117 22936
rect 52151 22933 52163 22967
rect 52105 22927 52163 22933
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 26605 22763 26663 22769
rect 26605 22729 26617 22763
rect 26651 22760 26663 22763
rect 27062 22760 27068 22772
rect 26651 22732 27068 22760
rect 26651 22729 26663 22732
rect 26605 22723 26663 22729
rect 27062 22720 27068 22732
rect 27120 22720 27126 22772
rect 28994 22760 29000 22772
rect 28955 22732 29000 22760
rect 28994 22720 29000 22732
rect 29052 22720 29058 22772
rect 37734 22720 37740 22772
rect 37792 22760 37798 22772
rect 37829 22763 37887 22769
rect 37829 22760 37841 22763
rect 37792 22732 37841 22760
rect 37792 22720 37798 22732
rect 37829 22729 37841 22732
rect 37875 22729 37887 22763
rect 37829 22723 37887 22729
rect 39393 22763 39451 22769
rect 39393 22729 39405 22763
rect 39439 22729 39451 22763
rect 40494 22760 40500 22772
rect 40455 22732 40500 22760
rect 39393 22723 39451 22729
rect 2406 22652 2412 22704
rect 2464 22692 2470 22704
rect 2464 22664 33350 22692
rect 2464 22652 2470 22664
rect 37274 22652 37280 22704
rect 37332 22692 37338 22704
rect 37645 22695 37703 22701
rect 37645 22692 37657 22695
rect 37332 22664 37657 22692
rect 37332 22652 37338 22664
rect 37645 22661 37657 22664
rect 37691 22661 37703 22695
rect 37645 22655 37703 22661
rect 39022 22652 39028 22704
rect 39080 22692 39086 22704
rect 39301 22695 39359 22701
rect 39301 22692 39313 22695
rect 39080 22664 39313 22692
rect 39080 22652 39086 22664
rect 39301 22661 39313 22664
rect 39347 22661 39359 22695
rect 39408 22692 39436 22723
rect 40494 22720 40500 22732
rect 40552 22720 40558 22772
rect 41690 22720 41696 22772
rect 41748 22760 41754 22772
rect 41969 22763 42027 22769
rect 41969 22760 41981 22763
rect 41748 22732 41981 22760
rect 41748 22720 41754 22732
rect 41969 22729 41981 22732
rect 42015 22760 42027 22763
rect 42426 22760 42432 22772
rect 42015 22732 42432 22760
rect 42015 22729 42027 22732
rect 41969 22723 42027 22729
rect 42426 22720 42432 22732
rect 42484 22760 42490 22772
rect 42484 22732 43300 22760
rect 42484 22720 42490 22732
rect 42886 22692 42892 22704
rect 39408 22664 40724 22692
rect 42847 22664 42892 22692
rect 39301 22655 39359 22661
rect 25961 22627 26019 22633
rect 25961 22593 25973 22627
rect 26007 22624 26019 22627
rect 26694 22624 26700 22636
rect 26007 22596 26700 22624
rect 26007 22593 26019 22596
rect 25961 22587 26019 22593
rect 26694 22584 26700 22596
rect 26752 22584 26758 22636
rect 28810 22584 28816 22636
rect 28868 22624 28874 22636
rect 29454 22624 29460 22636
rect 28868 22596 28913 22624
rect 29415 22596 29460 22624
rect 28868 22584 28874 22596
rect 29454 22584 29460 22596
rect 29512 22584 29518 22636
rect 29917 22627 29975 22633
rect 29917 22624 29929 22627
rect 29564 22596 29929 22624
rect 22830 22516 22836 22568
rect 22888 22556 22894 22568
rect 23569 22559 23627 22565
rect 23569 22556 23581 22559
rect 22888 22528 23581 22556
rect 22888 22516 22894 22528
rect 23569 22525 23581 22528
rect 23615 22525 23627 22559
rect 23569 22519 23627 22525
rect 26053 22559 26111 22565
rect 26053 22525 26065 22559
rect 26099 22556 26111 22559
rect 26234 22556 26240 22568
rect 26099 22528 26240 22556
rect 26099 22525 26111 22528
rect 26053 22519 26111 22525
rect 26234 22516 26240 22528
rect 26292 22556 26298 22568
rect 26970 22556 26976 22568
rect 26292 22528 26976 22556
rect 26292 22516 26298 22528
rect 26970 22516 26976 22528
rect 27028 22516 27034 22568
rect 27522 22516 27528 22568
rect 27580 22556 27586 22568
rect 28534 22556 28540 22568
rect 27580 22528 28540 22556
rect 27580 22516 27586 22528
rect 28534 22516 28540 22528
rect 28592 22516 28598 22568
rect 23293 22491 23351 22497
rect 23293 22457 23305 22491
rect 23339 22488 23351 22491
rect 23382 22488 23388 22500
rect 23339 22460 23388 22488
rect 23339 22457 23351 22460
rect 23293 22451 23351 22457
rect 23382 22448 23388 22460
rect 23440 22448 23446 22500
rect 25038 22448 25044 22500
rect 25096 22488 25102 22500
rect 28629 22491 28687 22497
rect 28629 22488 28641 22491
rect 25096 22460 28641 22488
rect 25096 22448 25102 22460
rect 28629 22457 28641 22460
rect 28675 22457 28687 22491
rect 28629 22451 28687 22457
rect 23106 22420 23112 22432
rect 23067 22392 23112 22420
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 24949 22423 25007 22429
rect 24949 22389 24961 22423
rect 24995 22420 25007 22423
rect 25866 22420 25872 22432
rect 24995 22392 25872 22420
rect 24995 22389 25007 22392
rect 24949 22383 25007 22389
rect 25866 22380 25872 22392
rect 25924 22380 25930 22432
rect 28644 22420 28672 22451
rect 29564 22420 29592 22596
rect 29917 22593 29929 22596
rect 29963 22593 29975 22627
rect 30282 22624 30288 22636
rect 30243 22596 30288 22624
rect 29917 22587 29975 22593
rect 30282 22584 30288 22596
rect 30340 22584 30346 22636
rect 30558 22584 30564 22636
rect 30616 22624 30622 22636
rect 30653 22627 30711 22633
rect 30653 22624 30665 22627
rect 30616 22596 30665 22624
rect 30616 22584 30622 22596
rect 30653 22593 30665 22596
rect 30699 22593 30711 22627
rect 31018 22624 31024 22636
rect 30979 22596 31024 22624
rect 30653 22587 30711 22593
rect 31018 22584 31024 22596
rect 31076 22584 31082 22636
rect 31294 22624 31300 22636
rect 31255 22596 31300 22624
rect 31294 22584 31300 22596
rect 31352 22624 31358 22636
rect 31846 22624 31852 22636
rect 31352 22596 31852 22624
rect 31352 22584 31358 22596
rect 31846 22584 31852 22596
rect 31904 22584 31910 22636
rect 33962 22624 33968 22636
rect 33923 22596 33968 22624
rect 33962 22584 33968 22596
rect 34020 22584 34026 22636
rect 34790 22624 34796 22636
rect 34751 22596 34796 22624
rect 34790 22584 34796 22596
rect 34848 22584 34854 22636
rect 37458 22624 37464 22636
rect 37419 22596 37464 22624
rect 37458 22584 37464 22596
rect 37516 22584 37522 22636
rect 39117 22627 39175 22633
rect 39117 22593 39129 22627
rect 39163 22624 39175 22627
rect 39206 22624 39212 22636
rect 39163 22596 39212 22624
rect 39163 22593 39175 22596
rect 39117 22587 39175 22593
rect 39206 22584 39212 22596
rect 39264 22584 39270 22636
rect 39868 22633 39896 22664
rect 39393 22627 39451 22633
rect 39393 22593 39405 22627
rect 39439 22593 39451 22627
rect 39393 22587 39451 22593
rect 39853 22627 39911 22633
rect 39853 22593 39865 22627
rect 39899 22593 39911 22627
rect 39853 22587 39911 22593
rect 39114 22448 39120 22500
rect 39172 22488 39178 22500
rect 39408 22488 39436 22587
rect 40126 22584 40132 22636
rect 40184 22624 40190 22636
rect 40494 22624 40500 22636
rect 40184 22596 40500 22624
rect 40184 22584 40190 22596
rect 40494 22584 40500 22596
rect 40552 22584 40558 22636
rect 40696 22633 40724 22664
rect 42886 22652 42892 22664
rect 42944 22652 42950 22704
rect 43272 22692 43300 22732
rect 44174 22720 44180 22772
rect 44232 22760 44238 22772
rect 44361 22763 44419 22769
rect 44361 22760 44373 22763
rect 44232 22732 44373 22760
rect 44232 22720 44238 22732
rect 44361 22729 44373 22732
rect 44407 22729 44419 22763
rect 44361 22723 44419 22729
rect 45925 22763 45983 22769
rect 45925 22729 45937 22763
rect 45971 22760 45983 22763
rect 46014 22760 46020 22772
rect 45971 22732 46020 22760
rect 45971 22729 45983 22732
rect 45925 22723 45983 22729
rect 46014 22720 46020 22732
rect 46072 22760 46078 22772
rect 46569 22763 46627 22769
rect 46569 22760 46581 22763
rect 46072 22732 46581 22760
rect 46072 22720 46078 22732
rect 46569 22729 46581 22732
rect 46615 22760 46627 22763
rect 46658 22760 46664 22772
rect 46615 22732 46664 22760
rect 46615 22729 46627 22732
rect 46569 22723 46627 22729
rect 46658 22720 46664 22732
rect 46716 22720 46722 22772
rect 47949 22763 48007 22769
rect 47949 22760 47961 22763
rect 46768 22732 47961 22760
rect 46768 22704 46796 22732
rect 47949 22729 47961 22732
rect 47995 22729 48007 22763
rect 47949 22723 48007 22729
rect 48038 22720 48044 22772
rect 48096 22760 48102 22772
rect 50985 22763 51043 22769
rect 48096 22732 48141 22760
rect 48096 22720 48102 22732
rect 50985 22729 50997 22763
rect 51031 22760 51043 22763
rect 51994 22760 52000 22772
rect 51031 22732 52000 22760
rect 51031 22729 51043 22732
rect 50985 22723 51043 22729
rect 51994 22720 52000 22732
rect 52052 22720 52058 22772
rect 56962 22760 56968 22772
rect 56923 22732 56968 22760
rect 56962 22720 56968 22732
rect 57020 22720 57026 22772
rect 58158 22760 58164 22772
rect 58119 22732 58164 22760
rect 58158 22720 58164 22732
rect 58216 22720 58222 22772
rect 45465 22695 45523 22701
rect 43272 22664 43378 22692
rect 45465 22661 45477 22695
rect 45511 22692 45523 22695
rect 46750 22692 46756 22704
rect 45511 22664 46756 22692
rect 45511 22661 45523 22664
rect 45465 22655 45523 22661
rect 46750 22652 46756 22664
rect 46808 22652 46814 22704
rect 47302 22652 47308 22704
rect 47360 22692 47366 22704
rect 48133 22695 48191 22701
rect 48133 22692 48145 22695
rect 47360 22664 48145 22692
rect 47360 22652 47366 22664
rect 48133 22661 48145 22664
rect 48179 22661 48191 22695
rect 54662 22692 54668 22704
rect 48133 22655 48191 22661
rect 54128 22664 54668 22692
rect 40681 22627 40739 22633
rect 40681 22593 40693 22627
rect 40727 22593 40739 22627
rect 40681 22587 40739 22593
rect 40770 22584 40776 22636
rect 40828 22624 40834 22636
rect 41141 22627 41199 22633
rect 41141 22624 41153 22627
rect 40828 22596 41153 22624
rect 40828 22584 40834 22596
rect 41141 22593 41153 22596
rect 41187 22593 41199 22627
rect 41322 22624 41328 22636
rect 41283 22596 41328 22624
rect 41141 22587 41199 22593
rect 41322 22584 41328 22596
rect 41380 22584 41386 22636
rect 45738 22624 45744 22636
rect 45651 22596 45744 22624
rect 45738 22584 45744 22596
rect 45796 22624 45802 22636
rect 46198 22624 46204 22636
rect 45796 22596 46204 22624
rect 45796 22584 45802 22596
rect 46198 22584 46204 22596
rect 46256 22584 46262 22636
rect 46566 22584 46572 22636
rect 46624 22624 46630 22636
rect 47765 22627 47823 22633
rect 47765 22624 47777 22627
rect 46624 22596 47777 22624
rect 46624 22584 46630 22596
rect 47765 22593 47777 22596
rect 47811 22593 47823 22627
rect 47765 22587 47823 22593
rect 49234 22584 49240 22636
rect 49292 22624 49298 22636
rect 49329 22627 49387 22633
rect 49329 22624 49341 22627
rect 49292 22596 49341 22624
rect 49292 22584 49298 22596
rect 49329 22593 49341 22596
rect 49375 22593 49387 22627
rect 49329 22587 49387 22593
rect 49513 22627 49571 22633
rect 49513 22593 49525 22627
rect 49559 22624 49571 22627
rect 50617 22627 50675 22633
rect 50617 22624 50629 22627
rect 49559 22596 50629 22624
rect 49559 22593 49571 22596
rect 49513 22587 49571 22593
rect 50617 22593 50629 22596
rect 50663 22624 50675 22627
rect 51258 22624 51264 22636
rect 50663 22596 51264 22624
rect 50663 22593 50675 22596
rect 50617 22587 50675 22593
rect 51258 22584 51264 22596
rect 51316 22584 51322 22636
rect 51718 22624 51724 22636
rect 51679 22596 51724 22624
rect 51718 22584 51724 22596
rect 51776 22584 51782 22636
rect 53374 22624 53380 22636
rect 53335 22596 53380 22624
rect 53374 22584 53380 22596
rect 53432 22584 53438 22636
rect 53558 22624 53564 22636
rect 53519 22596 53564 22624
rect 53558 22584 53564 22596
rect 53616 22584 53622 22636
rect 53742 22584 53748 22636
rect 53800 22624 53806 22636
rect 54128 22633 54156 22664
rect 54662 22652 54668 22664
rect 54720 22652 54726 22704
rect 56594 22692 56600 22704
rect 56555 22664 56600 22692
rect 56594 22652 56600 22664
rect 56652 22652 56658 22704
rect 56778 22652 56784 22704
rect 56836 22701 56842 22704
rect 56836 22695 56855 22701
rect 56843 22661 56855 22695
rect 56836 22655 56855 22661
rect 56836 22652 56842 22655
rect 53837 22627 53895 22633
rect 53837 22624 53849 22627
rect 53800 22596 53849 22624
rect 53800 22584 53806 22596
rect 53837 22593 53849 22596
rect 53883 22593 53895 22627
rect 53837 22587 53895 22593
rect 54113 22627 54171 22633
rect 54113 22593 54125 22627
rect 54159 22593 54171 22627
rect 54113 22587 54171 22593
rect 54205 22627 54263 22633
rect 54205 22593 54217 22627
rect 54251 22593 54263 22627
rect 54205 22587 54263 22593
rect 54941 22627 54999 22633
rect 54941 22593 54953 22627
rect 54987 22593 54999 22627
rect 55122 22624 55128 22636
rect 55083 22596 55128 22624
rect 54941 22587 54999 22593
rect 39945 22559 40003 22565
rect 39945 22525 39957 22559
rect 39991 22556 40003 22559
rect 40586 22556 40592 22568
rect 39991 22528 40592 22556
rect 39991 22525 40003 22528
rect 39945 22519 40003 22525
rect 40586 22516 40592 22528
rect 40644 22516 40650 22568
rect 41598 22516 41604 22568
rect 41656 22556 41662 22568
rect 42613 22559 42671 22565
rect 42613 22556 42625 22559
rect 41656 22528 42625 22556
rect 41656 22516 41662 22528
rect 42613 22525 42625 22528
rect 42659 22525 42671 22559
rect 45646 22556 45652 22568
rect 45607 22528 45652 22556
rect 42613 22519 42671 22525
rect 39172 22460 39436 22488
rect 39172 22448 39178 22460
rect 28644 22392 29592 22420
rect 41233 22423 41291 22429
rect 41233 22389 41245 22423
rect 41279 22420 41291 22423
rect 41506 22420 41512 22432
rect 41279 22392 41512 22420
rect 41279 22389 41291 22392
rect 41233 22383 41291 22389
rect 41506 22380 41512 22392
rect 41564 22380 41570 22432
rect 42628 22420 42656 22519
rect 45646 22516 45652 22528
rect 45704 22516 45710 22568
rect 46017 22559 46075 22565
rect 46017 22525 46029 22559
rect 46063 22525 46075 22559
rect 46017 22519 46075 22525
rect 44913 22491 44971 22497
rect 44913 22457 44925 22491
rect 44959 22488 44971 22491
rect 45554 22488 45560 22500
rect 44959 22460 45560 22488
rect 44959 22457 44971 22460
rect 44913 22451 44971 22457
rect 44928 22420 44956 22451
rect 45554 22448 45560 22460
rect 45612 22448 45618 22500
rect 42628 22392 44956 22420
rect 46032 22420 46060 22519
rect 46106 22516 46112 22568
rect 46164 22556 46170 22568
rect 46164 22528 46209 22556
rect 46164 22516 46170 22528
rect 49694 22516 49700 22568
rect 49752 22556 49758 22568
rect 50525 22559 50583 22565
rect 50525 22556 50537 22559
rect 49752 22528 50537 22556
rect 49752 22516 49758 22528
rect 50525 22525 50537 22528
rect 50571 22525 50583 22559
rect 50525 22519 50583 22525
rect 51629 22559 51687 22565
rect 51629 22525 51641 22559
rect 51675 22525 51687 22559
rect 52086 22556 52092 22568
rect 52047 22528 52092 22556
rect 51629 22519 51687 22525
rect 48317 22491 48375 22497
rect 48317 22457 48329 22491
rect 48363 22488 48375 22491
rect 51644 22488 51672 22519
rect 52086 22516 52092 22528
rect 52144 22516 52150 22568
rect 52178 22516 52184 22568
rect 52236 22556 52242 22568
rect 53650 22556 53656 22568
rect 52236 22528 53656 22556
rect 52236 22516 52242 22528
rect 53650 22516 53656 22528
rect 53708 22556 53714 22568
rect 54220 22556 54248 22587
rect 53708 22528 54248 22556
rect 54956 22556 54984 22587
rect 55122 22584 55128 22596
rect 55180 22584 55186 22636
rect 55582 22624 55588 22636
rect 55543 22596 55588 22624
rect 55582 22584 55588 22596
rect 55640 22584 55646 22636
rect 55858 22556 55864 22568
rect 54956 22528 55864 22556
rect 53708 22516 53714 22528
rect 55858 22516 55864 22528
rect 55916 22516 55922 22568
rect 52638 22488 52644 22500
rect 48363 22460 52644 22488
rect 48363 22457 48375 22460
rect 48317 22451 48375 22457
rect 52638 22448 52644 22460
rect 52696 22448 52702 22500
rect 47213 22423 47271 22429
rect 47213 22420 47225 22423
rect 46032 22392 47225 22420
rect 47213 22389 47225 22392
rect 47259 22420 47271 22423
rect 47670 22420 47676 22432
rect 47259 22392 47676 22420
rect 47259 22389 47271 22392
rect 47213 22383 47271 22389
rect 47670 22380 47676 22392
rect 47728 22380 47734 22432
rect 49418 22380 49424 22432
rect 49476 22420 49482 22432
rect 49513 22423 49571 22429
rect 49513 22420 49525 22423
rect 49476 22392 49525 22420
rect 49476 22380 49482 22392
rect 49513 22389 49525 22392
rect 49559 22389 49571 22423
rect 49513 22383 49571 22389
rect 55033 22423 55091 22429
rect 55033 22389 55045 22423
rect 55079 22420 55091 22423
rect 55674 22420 55680 22432
rect 55079 22392 55680 22420
rect 55079 22389 55091 22392
rect 55033 22383 55091 22389
rect 55674 22380 55680 22392
rect 55732 22380 55738 22432
rect 56045 22423 56103 22429
rect 56045 22389 56057 22423
rect 56091 22420 56103 22423
rect 56502 22420 56508 22432
rect 56091 22392 56508 22420
rect 56091 22389 56103 22392
rect 56045 22383 56103 22389
rect 56502 22380 56508 22392
rect 56560 22420 56566 22432
rect 56781 22423 56839 22429
rect 56781 22420 56793 22423
rect 56560 22392 56793 22420
rect 56560 22380 56566 22392
rect 56781 22389 56793 22392
rect 56827 22389 56839 22423
rect 56781 22383 56839 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 27522 22216 27528 22228
rect 27483 22188 27528 22216
rect 27522 22176 27528 22188
rect 27580 22176 27586 22228
rect 27985 22219 28043 22225
rect 27985 22185 27997 22219
rect 28031 22185 28043 22219
rect 27985 22179 28043 22185
rect 28353 22219 28411 22225
rect 28353 22185 28365 22219
rect 28399 22216 28411 22219
rect 28626 22216 28632 22228
rect 28399 22188 28632 22216
rect 28399 22185 28411 22188
rect 28353 22179 28411 22185
rect 24762 22080 24768 22092
rect 23952 22052 24768 22080
rect 23106 21972 23112 22024
rect 23164 22012 23170 22024
rect 23382 22012 23388 22024
rect 23164 21984 23388 22012
rect 23164 21972 23170 21984
rect 23382 21972 23388 21984
rect 23440 22012 23446 22024
rect 23952 22021 23980 22052
rect 24762 22040 24768 22052
rect 24820 22040 24826 22092
rect 25038 22080 25044 22092
rect 24999 22052 25044 22080
rect 25038 22040 25044 22052
rect 25096 22040 25102 22092
rect 28000 22080 28028 22179
rect 28626 22176 28632 22188
rect 28684 22176 28690 22228
rect 30742 22216 30748 22228
rect 30703 22188 30748 22216
rect 30742 22176 30748 22188
rect 30800 22176 30806 22228
rect 34790 22216 34796 22228
rect 31772 22188 34796 22216
rect 31772 22080 31800 22188
rect 34790 22176 34796 22188
rect 34848 22216 34854 22228
rect 34885 22219 34943 22225
rect 34885 22216 34897 22219
rect 34848 22188 34897 22216
rect 34848 22176 34854 22188
rect 34885 22185 34897 22188
rect 34931 22185 34943 22219
rect 34885 22179 34943 22185
rect 42426 22176 42432 22228
rect 42484 22216 42490 22228
rect 42705 22219 42763 22225
rect 42705 22216 42717 22219
rect 42484 22188 42717 22216
rect 42484 22176 42490 22188
rect 42705 22185 42717 22188
rect 42751 22185 42763 22219
rect 42705 22179 42763 22185
rect 44358 22176 44364 22228
rect 44416 22216 44422 22228
rect 44453 22219 44511 22225
rect 44453 22216 44465 22219
rect 44416 22188 44465 22216
rect 44416 22176 44422 22188
rect 44453 22185 44465 22188
rect 44499 22185 44511 22219
rect 44453 22179 44511 22185
rect 44542 22176 44548 22228
rect 44600 22216 44606 22228
rect 48869 22219 48927 22225
rect 44600 22188 46888 22216
rect 44600 22176 44606 22188
rect 32582 22108 32588 22160
rect 32640 22148 32646 22160
rect 33321 22151 33379 22157
rect 33321 22148 33333 22151
rect 32640 22120 33333 22148
rect 32640 22108 32646 22120
rect 33321 22117 33333 22120
rect 33367 22117 33379 22151
rect 43625 22151 43683 22157
rect 33321 22111 33379 22117
rect 40972 22120 41828 22148
rect 40972 22092 41000 22120
rect 27172 22052 28028 22080
rect 31680 22052 31800 22080
rect 27172 22024 27200 22052
rect 23937 22015 23995 22021
rect 23440 21984 23888 22012
rect 23440 21972 23446 21984
rect 23750 21944 23756 21956
rect 23711 21916 23756 21944
rect 23750 21904 23756 21916
rect 23808 21904 23814 21956
rect 23860 21944 23888 21984
rect 23937 21981 23949 22015
rect 23983 21981 23995 22015
rect 23937 21975 23995 21981
rect 24026 21972 24032 22024
rect 24084 22012 24090 22024
rect 24084 21984 24129 22012
rect 24084 21972 24090 21984
rect 24670 21972 24676 22024
rect 24728 22012 24734 22024
rect 24857 22015 24915 22021
rect 24857 22012 24869 22015
rect 24728 21984 24869 22012
rect 24728 21972 24734 21984
rect 24857 21981 24869 21984
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 25682 21972 25688 22024
rect 25740 22012 25746 22024
rect 25866 22012 25872 22024
rect 25740 21984 25872 22012
rect 25740 21972 25746 21984
rect 25866 21972 25872 21984
rect 25924 22012 25930 22024
rect 25961 22015 26019 22021
rect 25961 22012 25973 22015
rect 25924 21984 25973 22012
rect 25924 21972 25930 21984
rect 25961 21981 25973 21984
rect 26007 21981 26019 22015
rect 25961 21975 26019 21981
rect 26329 22015 26387 22021
rect 26329 21981 26341 22015
rect 26375 22012 26387 22015
rect 26418 22012 26424 22024
rect 26375 21984 26424 22012
rect 26375 21981 26387 21984
rect 26329 21975 26387 21981
rect 26418 21972 26424 21984
rect 26476 21972 26482 22024
rect 27062 22012 27068 22024
rect 27023 21984 27068 22012
rect 27062 21972 27068 21984
rect 27120 21972 27126 22024
rect 27154 21972 27160 22024
rect 27212 22012 27218 22024
rect 27341 22015 27399 22021
rect 27212 21984 27257 22012
rect 27212 21972 27218 21984
rect 27341 21981 27353 22015
rect 27387 22012 27399 22015
rect 27706 22012 27712 22024
rect 27387 21984 27712 22012
rect 27387 21981 27399 21984
rect 27341 21975 27399 21981
rect 27706 21972 27712 21984
rect 27764 22012 27770 22024
rect 27985 22015 28043 22021
rect 27985 22012 27997 22015
rect 27764 21984 27997 22012
rect 27764 21972 27770 21984
rect 27985 21981 27997 21984
rect 28031 21981 28043 22015
rect 27985 21975 28043 21981
rect 28077 22015 28135 22021
rect 28077 21981 28089 22015
rect 28123 21981 28135 22015
rect 28077 21975 28135 21981
rect 30929 22015 30987 22021
rect 30929 21981 30941 22015
rect 30975 21981 30987 22015
rect 31110 22012 31116 22024
rect 31071 21984 31116 22012
rect 30929 21975 30987 21981
rect 24581 21947 24639 21953
rect 24581 21944 24593 21947
rect 23860 21916 24593 21944
rect 24581 21913 24593 21916
rect 24627 21913 24639 21947
rect 27080 21944 27108 21972
rect 28092 21944 28120 21975
rect 27080 21916 28120 21944
rect 30944 21944 30972 21975
rect 31110 21972 31116 21984
rect 31168 21972 31174 22024
rect 31205 22015 31263 22021
rect 31205 21981 31217 22015
rect 31251 22012 31263 22015
rect 31294 22012 31300 22024
rect 31251 21984 31300 22012
rect 31251 21981 31263 21984
rect 31205 21975 31263 21981
rect 31294 21972 31300 21984
rect 31352 21972 31358 22024
rect 31680 22021 31708 22052
rect 31846 22040 31852 22092
rect 31904 22080 31910 22092
rect 33781 22083 33839 22089
rect 31904 22052 32076 22080
rect 31904 22040 31910 22052
rect 31665 22015 31723 22021
rect 31665 21981 31677 22015
rect 31711 21981 31723 22015
rect 31665 21975 31723 21981
rect 31754 21972 31760 22024
rect 31812 22012 31818 22024
rect 32048 22021 32076 22052
rect 33781 22049 33793 22083
rect 33827 22080 33839 22083
rect 34514 22080 34520 22092
rect 33827 22052 34520 22080
rect 33827 22049 33839 22052
rect 33781 22043 33839 22049
rect 34514 22040 34520 22052
rect 34572 22040 34578 22092
rect 38930 22040 38936 22092
rect 38988 22080 38994 22092
rect 39485 22083 39543 22089
rect 38988 22052 39436 22080
rect 38988 22040 38994 22052
rect 32033 22015 32091 22021
rect 31812 21984 31857 22012
rect 31812 21972 31818 21984
rect 32033 21981 32045 22015
rect 32079 21981 32091 22015
rect 32033 21975 32091 21981
rect 32122 21972 32128 22024
rect 32180 22012 32186 22024
rect 32180 21984 32225 22012
rect 32180 21972 32186 21984
rect 33318 21972 33324 22024
rect 33376 22012 33382 22024
rect 33689 22015 33747 22021
rect 33689 22012 33701 22015
rect 33376 21984 33701 22012
rect 33376 21972 33382 21984
rect 33689 21981 33701 21984
rect 33735 21981 33747 22015
rect 35526 22012 35532 22024
rect 35487 21984 35532 22012
rect 33689 21975 33747 21981
rect 35526 21972 35532 21984
rect 35584 21972 35590 22024
rect 36357 22015 36415 22021
rect 36357 21981 36369 22015
rect 36403 21981 36415 22015
rect 39022 22012 39028 22024
rect 38983 21984 39028 22012
rect 36357 21975 36415 21981
rect 31938 21944 31944 21956
rect 30944 21916 31754 21944
rect 31899 21916 31944 21944
rect 24581 21907 24639 21913
rect 31726 21888 31754 21916
rect 31938 21904 31944 21916
rect 31996 21904 32002 21956
rect 35434 21904 35440 21956
rect 35492 21944 35498 21956
rect 36372 21944 36400 21975
rect 39022 21972 39028 21984
rect 39080 21972 39086 22024
rect 39298 22012 39304 22024
rect 39259 21984 39304 22012
rect 39298 21972 39304 21984
rect 39356 21972 39362 22024
rect 39408 22012 39436 22052
rect 39485 22049 39497 22083
rect 39531 22080 39543 22083
rect 40494 22080 40500 22092
rect 39531 22052 40500 22080
rect 39531 22049 39543 22052
rect 39485 22043 39543 22049
rect 40494 22040 40500 22052
rect 40552 22040 40558 22092
rect 40770 22080 40776 22092
rect 40604 22052 40776 22080
rect 40604 22012 40632 22052
rect 40770 22040 40776 22052
rect 40828 22040 40834 22092
rect 40954 22040 40960 22092
rect 41012 22040 41018 22092
rect 41800 22080 41828 22120
rect 43625 22117 43637 22151
rect 43671 22148 43683 22151
rect 45554 22148 45560 22160
rect 43671 22120 45560 22148
rect 43671 22117 43683 22120
rect 43625 22111 43683 22117
rect 45554 22108 45560 22120
rect 45612 22108 45618 22160
rect 46290 22108 46296 22160
rect 46348 22148 46354 22160
rect 46753 22151 46811 22157
rect 46753 22148 46765 22151
rect 46348 22120 46765 22148
rect 46348 22108 46354 22120
rect 46753 22117 46765 22120
rect 46799 22117 46811 22151
rect 46860 22148 46888 22188
rect 48869 22185 48881 22219
rect 48915 22216 48927 22219
rect 48958 22216 48964 22228
rect 48915 22188 48964 22216
rect 48915 22185 48927 22188
rect 48869 22179 48927 22185
rect 48958 22176 48964 22188
rect 49016 22176 49022 22228
rect 50801 22219 50859 22225
rect 50801 22185 50813 22219
rect 50847 22216 50859 22219
rect 53098 22216 53104 22228
rect 50847 22188 53104 22216
rect 50847 22185 50859 22188
rect 50801 22179 50859 22185
rect 53098 22176 53104 22188
rect 53156 22176 53162 22228
rect 53282 22216 53288 22228
rect 53243 22188 53288 22216
rect 53282 22176 53288 22188
rect 53340 22176 53346 22228
rect 56781 22219 56839 22225
rect 56781 22185 56793 22219
rect 56827 22216 56839 22219
rect 57422 22216 57428 22228
rect 56827 22188 57428 22216
rect 56827 22185 56839 22188
rect 56781 22179 56839 22185
rect 57422 22176 57428 22188
rect 57480 22176 57486 22228
rect 58066 22176 58072 22228
rect 58124 22216 58130 22228
rect 58161 22219 58219 22225
rect 58161 22216 58173 22219
rect 58124 22188 58173 22216
rect 58124 22176 58130 22188
rect 58161 22185 58173 22188
rect 58207 22185 58219 22219
rect 58161 22179 58219 22185
rect 57974 22148 57980 22160
rect 46860 22120 57980 22148
rect 46753 22111 46811 22117
rect 57974 22108 57980 22120
rect 58032 22108 58038 22160
rect 41969 22083 42027 22089
rect 41969 22080 41981 22083
rect 41064 22052 41414 22080
rect 41800 22052 41981 22080
rect 39408 21984 40632 22012
rect 40681 22015 40739 22021
rect 40681 21981 40693 22015
rect 40727 22012 40739 22015
rect 40972 22012 41000 22040
rect 41064 22021 41092 22052
rect 40727 21984 41000 22012
rect 41049 22015 41107 22021
rect 40727 21981 40739 21984
rect 40681 21975 40739 21981
rect 41049 21981 41061 22015
rect 41095 21981 41107 22015
rect 41049 21975 41107 21981
rect 41138 21972 41144 22024
rect 41196 22012 41202 22024
rect 41386 22012 41414 22052
rect 41969 22049 41981 22052
rect 42015 22049 42027 22083
rect 41969 22043 42027 22049
rect 47213 22083 47271 22089
rect 47213 22049 47225 22083
rect 47259 22080 47271 22083
rect 47762 22080 47768 22092
rect 47259 22052 47768 22080
rect 47259 22049 47271 22052
rect 47213 22043 47271 22049
rect 47762 22040 47768 22052
rect 47820 22040 47826 22092
rect 47854 22040 47860 22092
rect 47912 22080 47918 22092
rect 49234 22080 49240 22092
rect 47912 22052 49240 22080
rect 47912 22040 47918 22052
rect 49234 22040 49240 22052
rect 49292 22040 49298 22092
rect 49329 22083 49387 22089
rect 49329 22049 49341 22083
rect 49375 22080 49387 22083
rect 49418 22080 49424 22092
rect 49375 22052 49424 22080
rect 49375 22049 49387 22052
rect 49329 22043 49387 22049
rect 49418 22040 49424 22052
rect 49476 22040 49482 22092
rect 50154 22040 50160 22092
rect 50212 22080 50218 22092
rect 50433 22083 50491 22089
rect 50433 22080 50445 22083
rect 50212 22052 50445 22080
rect 50212 22040 50218 22052
rect 50433 22049 50445 22052
rect 50479 22049 50491 22083
rect 53558 22080 53564 22092
rect 53471 22052 53564 22080
rect 50433 22043 50491 22049
rect 53558 22040 53564 22052
rect 53616 22080 53622 22092
rect 54389 22083 54447 22089
rect 54389 22080 54401 22083
rect 53616 22052 54401 22080
rect 53616 22040 53622 22052
rect 54389 22049 54401 22052
rect 54435 22049 54447 22083
rect 55858 22080 55864 22092
rect 55819 22052 55864 22080
rect 54389 22043 54447 22049
rect 55858 22040 55864 22052
rect 55916 22040 55922 22092
rect 57790 22080 57796 22092
rect 57751 22052 57796 22080
rect 57790 22040 57796 22052
rect 57848 22040 57854 22092
rect 41690 22012 41696 22024
rect 41196 21984 41241 22012
rect 41386 21984 41696 22012
rect 41196 21972 41202 21984
rect 41690 21972 41696 21984
rect 41748 21972 41754 22024
rect 41785 22015 41843 22021
rect 41785 21981 41797 22015
rect 41831 21981 41843 22015
rect 41785 21975 41843 21981
rect 41877 22015 41935 22021
rect 41877 21981 41889 22015
rect 41923 21981 41935 22015
rect 41877 21975 41935 21981
rect 44177 22015 44235 22021
rect 44177 21981 44189 22015
rect 44223 22012 44235 22015
rect 44818 22012 44824 22024
rect 44223 21984 44824 22012
rect 44223 21981 44235 21984
rect 44177 21975 44235 21981
rect 40770 21944 40776 21956
rect 35492 21916 40632 21944
rect 40731 21916 40776 21944
rect 35492 21904 35498 21916
rect 23842 21876 23848 21888
rect 23900 21885 23906 21888
rect 23809 21848 23848 21876
rect 23842 21836 23848 21848
rect 23900 21839 23909 21885
rect 23900 21836 23906 21839
rect 24486 21836 24492 21888
rect 24544 21876 24550 21888
rect 24673 21879 24731 21885
rect 24673 21876 24685 21879
rect 24544 21848 24685 21876
rect 24544 21836 24550 21848
rect 24673 21845 24685 21848
rect 24719 21845 24731 21879
rect 24673 21839 24731 21845
rect 24854 21836 24860 21888
rect 24912 21876 24918 21888
rect 25961 21879 26019 21885
rect 25961 21876 25973 21879
rect 24912 21848 25973 21876
rect 24912 21836 24918 21848
rect 25961 21845 25973 21848
rect 26007 21845 26019 21879
rect 25961 21839 26019 21845
rect 26050 21836 26056 21888
rect 26108 21876 26114 21888
rect 26145 21879 26203 21885
rect 26145 21876 26157 21879
rect 26108 21848 26157 21876
rect 26108 21836 26114 21848
rect 26145 21845 26157 21848
rect 26191 21845 26203 21879
rect 26145 21839 26203 21845
rect 26234 21836 26240 21888
rect 26292 21876 26298 21888
rect 26292 21848 26337 21876
rect 31726 21848 31760 21888
rect 26292 21836 26298 21848
rect 31754 21836 31760 21848
rect 31812 21836 31818 21888
rect 32309 21879 32367 21885
rect 32309 21845 32321 21879
rect 32355 21876 32367 21879
rect 38930 21876 38936 21888
rect 32355 21848 38936 21876
rect 32355 21845 32367 21848
rect 32309 21839 32367 21845
rect 38930 21836 38936 21848
rect 38988 21836 38994 21888
rect 39114 21876 39120 21888
rect 39075 21848 39120 21876
rect 39114 21836 39120 21848
rect 39172 21836 39178 21888
rect 40218 21836 40224 21888
rect 40276 21876 40282 21888
rect 40497 21879 40555 21885
rect 40497 21876 40509 21879
rect 40276 21848 40509 21876
rect 40276 21836 40282 21848
rect 40497 21845 40509 21848
rect 40543 21845 40555 21879
rect 40604 21876 40632 21916
rect 40770 21904 40776 21916
rect 40828 21904 40834 21956
rect 40862 21904 40868 21956
rect 40920 21944 40926 21956
rect 41322 21944 41328 21956
rect 40920 21916 41328 21944
rect 40920 21904 40926 21916
rect 41322 21904 41328 21916
rect 41380 21944 41386 21956
rect 41800 21944 41828 21975
rect 41380 21916 41828 21944
rect 41380 21904 41386 21916
rect 40678 21876 40684 21888
rect 40604 21848 40684 21876
rect 40497 21839 40555 21845
rect 40678 21836 40684 21848
rect 40736 21836 40742 21888
rect 40788 21876 40816 21904
rect 41892 21876 41920 21975
rect 44818 21972 44824 21984
rect 44876 21972 44882 22024
rect 45738 21972 45744 22024
rect 45796 22012 45802 22024
rect 45833 22015 45891 22021
rect 45833 22012 45845 22015
rect 45796 21984 45845 22012
rect 45796 21972 45802 21984
rect 45833 21981 45845 21984
rect 45879 21981 45891 22015
rect 47118 22012 47124 22024
rect 47079 21984 47124 22012
rect 45833 21975 45891 21981
rect 47118 21972 47124 21984
rect 47176 21972 47182 22024
rect 48774 21972 48780 22024
rect 48832 22012 48838 22024
rect 49053 22015 49111 22021
rect 49053 22012 49065 22015
rect 48832 21984 49065 22012
rect 48832 21972 48838 21984
rect 49053 21981 49065 21984
rect 49099 21981 49111 22015
rect 49053 21975 49111 21981
rect 49142 21972 49148 22024
rect 49200 22012 49206 22024
rect 49200 21984 49245 22012
rect 49200 21972 49206 21984
rect 50062 21972 50068 22024
rect 50120 22012 50126 22024
rect 50525 22015 50583 22021
rect 50525 22012 50537 22015
rect 50120 21984 50537 22012
rect 50120 21972 50126 21984
rect 50525 21981 50537 21984
rect 50571 21981 50583 22015
rect 50525 21975 50583 21981
rect 52457 22015 52515 22021
rect 52457 21981 52469 22015
rect 52503 22012 52515 22015
rect 53374 22012 53380 22024
rect 52503 21984 53380 22012
rect 52503 21981 52515 21984
rect 52457 21975 52515 21981
rect 53374 21972 53380 21984
rect 53432 22012 53438 22024
rect 53469 22015 53527 22021
rect 53469 22012 53481 22015
rect 53432 21984 53481 22012
rect 53432 21972 53438 21984
rect 53469 21981 53481 21984
rect 53515 21981 53527 22015
rect 53650 22012 53656 22024
rect 53611 21984 53656 22012
rect 53469 21975 53527 21981
rect 53650 21972 53656 21984
rect 53708 21972 53714 22024
rect 53742 21972 53748 22024
rect 53800 22012 53806 22024
rect 54297 22015 54355 22021
rect 53800 21984 53845 22012
rect 53800 21972 53806 21984
rect 54297 21981 54309 22015
rect 54343 22012 54355 22015
rect 54481 22015 54539 22021
rect 54343 21984 54432 22012
rect 54343 21981 54355 21984
rect 54297 21975 54355 21981
rect 44450 21944 44456 21956
rect 44411 21916 44456 21944
rect 44450 21904 44456 21916
rect 44508 21904 44514 21956
rect 52638 21944 52644 21956
rect 52599 21916 52644 21944
rect 52638 21904 52644 21916
rect 52696 21904 52702 21956
rect 52822 21944 52828 21956
rect 52783 21916 52828 21944
rect 52822 21904 52828 21916
rect 52880 21904 52886 21956
rect 53098 21904 53104 21956
rect 53156 21944 53162 21956
rect 53760 21944 53788 21972
rect 54404 21956 54432 21984
rect 54481 21981 54493 22015
rect 54527 21981 54539 22015
rect 54481 21975 54539 21981
rect 53156 21916 53788 21944
rect 53156 21904 53162 21916
rect 54386 21904 54392 21956
rect 54444 21904 54450 21956
rect 42150 21876 42156 21888
rect 40788 21848 41920 21876
rect 42111 21848 42156 21876
rect 42150 21836 42156 21848
rect 42208 21836 42214 21888
rect 44269 21879 44327 21885
rect 44269 21845 44281 21879
rect 44315 21876 44327 21879
rect 44910 21876 44916 21888
rect 44315 21848 44916 21876
rect 44315 21845 44327 21848
rect 44269 21839 44327 21845
rect 44910 21836 44916 21848
rect 44968 21876 44974 21888
rect 45370 21876 45376 21888
rect 44968 21848 45376 21876
rect 44968 21836 44974 21848
rect 45370 21836 45376 21848
rect 45428 21836 45434 21888
rect 46017 21879 46075 21885
rect 46017 21845 46029 21879
rect 46063 21876 46075 21879
rect 46566 21876 46572 21888
rect 46063 21848 46572 21876
rect 46063 21845 46075 21848
rect 46017 21839 46075 21845
rect 46566 21836 46572 21848
rect 46624 21836 46630 21888
rect 52656 21876 52684 21904
rect 54294 21876 54300 21888
rect 52656 21848 54300 21876
rect 54294 21836 54300 21848
rect 54352 21876 54358 21888
rect 54496 21876 54524 21975
rect 55214 21972 55220 22024
rect 55272 22012 55278 22024
rect 55677 22015 55735 22021
rect 55677 22012 55689 22015
rect 55272 21984 55689 22012
rect 55272 21972 55278 21984
rect 55677 21981 55689 21984
rect 55723 21981 55735 22015
rect 56502 22012 56508 22024
rect 56463 21984 56508 22012
rect 55677 21975 55735 21981
rect 56502 21972 56508 21984
rect 56560 21972 56566 22024
rect 57885 22015 57943 22021
rect 57885 21981 57897 22015
rect 57931 22012 57943 22015
rect 58158 22012 58164 22024
rect 57931 21984 58164 22012
rect 57931 21981 57943 21984
rect 57885 21975 57943 21981
rect 58158 21972 58164 21984
rect 58216 21972 58222 22024
rect 55030 21904 55036 21956
rect 55088 21944 55094 21956
rect 55493 21947 55551 21953
rect 55493 21944 55505 21947
rect 55088 21916 55505 21944
rect 55088 21904 55094 21916
rect 55493 21913 55505 21916
rect 55539 21913 55551 21947
rect 56778 21944 56784 21956
rect 56739 21916 56784 21944
rect 55493 21907 55551 21913
rect 56778 21904 56784 21916
rect 56836 21904 56842 21956
rect 54352 21848 54524 21876
rect 54352 21836 54358 21848
rect 55122 21836 55128 21888
rect 55180 21876 55186 21888
rect 56594 21876 56600 21888
rect 55180 21848 56600 21876
rect 55180 21836 55186 21848
rect 56594 21836 56600 21848
rect 56652 21836 56658 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 24486 21672 24492 21684
rect 24447 21644 24492 21672
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 24854 21672 24860 21684
rect 24815 21644 24860 21672
rect 24854 21632 24860 21644
rect 24912 21632 24918 21684
rect 26234 21632 26240 21684
rect 26292 21672 26298 21684
rect 26329 21675 26387 21681
rect 26329 21672 26341 21675
rect 26292 21644 26341 21672
rect 26292 21632 26298 21644
rect 26329 21641 26341 21644
rect 26375 21641 26387 21675
rect 26329 21635 26387 21641
rect 26605 21675 26663 21681
rect 26605 21641 26617 21675
rect 26651 21672 26663 21675
rect 27154 21672 27160 21684
rect 26651 21644 27160 21672
rect 26651 21641 26663 21644
rect 26605 21635 26663 21641
rect 27154 21632 27160 21644
rect 27212 21632 27218 21684
rect 27706 21672 27712 21684
rect 27667 21644 27712 21672
rect 27706 21632 27712 21644
rect 27764 21632 27770 21684
rect 31662 21632 31668 21684
rect 31720 21672 31726 21684
rect 31757 21675 31815 21681
rect 31757 21672 31769 21675
rect 31720 21644 31769 21672
rect 31720 21632 31726 21644
rect 31757 21641 31769 21644
rect 31803 21641 31815 21675
rect 31757 21635 31815 21641
rect 32122 21632 32128 21684
rect 32180 21672 32186 21684
rect 32585 21675 32643 21681
rect 32585 21672 32597 21675
rect 32180 21644 32597 21672
rect 32180 21632 32186 21644
rect 32585 21641 32597 21644
rect 32631 21641 32643 21675
rect 32585 21635 32643 21641
rect 36633 21675 36691 21681
rect 36633 21641 36645 21675
rect 36679 21672 36691 21675
rect 36722 21672 36728 21684
rect 36679 21644 36728 21672
rect 36679 21641 36691 21644
rect 36633 21635 36691 21641
rect 36722 21632 36728 21644
rect 36780 21632 36786 21684
rect 39025 21675 39083 21681
rect 39025 21641 39037 21675
rect 39071 21672 39083 21675
rect 39298 21672 39304 21684
rect 39071 21644 39304 21672
rect 39071 21641 39083 21644
rect 39025 21635 39083 21641
rect 39298 21632 39304 21644
rect 39356 21632 39362 21684
rect 40589 21675 40647 21681
rect 40589 21641 40601 21675
rect 40635 21672 40647 21675
rect 40862 21672 40868 21684
rect 40635 21644 40868 21672
rect 40635 21641 40647 21644
rect 40589 21635 40647 21641
rect 40862 21632 40868 21644
rect 40920 21632 40926 21684
rect 41230 21672 41236 21684
rect 41191 21644 41236 21672
rect 41230 21632 41236 21644
rect 41288 21632 41294 21684
rect 47762 21672 47768 21684
rect 47723 21644 47768 21672
rect 47762 21632 47768 21644
rect 47820 21632 47826 21684
rect 48774 21672 48780 21684
rect 48735 21644 48780 21672
rect 48774 21632 48780 21644
rect 48832 21632 48838 21684
rect 49234 21632 49240 21684
rect 49292 21672 49298 21684
rect 50062 21672 50068 21684
rect 49292 21644 50068 21672
rect 49292 21632 49298 21644
rect 50062 21632 50068 21644
rect 50120 21632 50126 21684
rect 52822 21632 52828 21684
rect 52880 21672 52886 21684
rect 54386 21672 54392 21684
rect 52880 21644 54392 21672
rect 52880 21632 52886 21644
rect 54386 21632 54392 21644
rect 54444 21632 54450 21684
rect 55122 21672 55128 21684
rect 55083 21644 55128 21672
rect 55122 21632 55128 21644
rect 55180 21632 55186 21684
rect 56778 21632 56784 21684
rect 56836 21672 56842 21684
rect 56965 21675 57023 21681
rect 56965 21672 56977 21675
rect 56836 21644 56977 21672
rect 56836 21632 56842 21644
rect 56965 21641 56977 21644
rect 57011 21641 57023 21675
rect 58158 21672 58164 21684
rect 58119 21644 58164 21672
rect 56965 21635 57023 21641
rect 58158 21632 58164 21644
rect 58216 21632 58222 21684
rect 24026 21564 24032 21616
rect 24084 21604 24090 21616
rect 27430 21604 27436 21616
rect 24084 21576 24992 21604
rect 24084 21564 24090 21576
rect 24964 21548 24992 21576
rect 25608 21576 27436 21604
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21536 23351 21539
rect 23658 21536 23664 21548
rect 23339 21508 23664 21536
rect 23339 21505 23351 21508
rect 23293 21499 23351 21505
rect 23658 21496 23664 21508
rect 23716 21496 23722 21548
rect 23750 21496 23756 21548
rect 23808 21536 23814 21548
rect 24673 21539 24731 21545
rect 24673 21536 24685 21539
rect 23808 21508 24685 21536
rect 23808 21496 23814 21508
rect 24673 21505 24685 21508
rect 24719 21536 24731 21539
rect 24762 21536 24768 21548
rect 24719 21508 24768 21536
rect 24719 21505 24731 21508
rect 24673 21499 24731 21505
rect 24762 21496 24768 21508
rect 24820 21496 24826 21548
rect 24946 21536 24952 21548
rect 24907 21508 24952 21536
rect 24946 21496 24952 21508
rect 25004 21496 25010 21548
rect 25038 21496 25044 21548
rect 25096 21536 25102 21548
rect 25608 21545 25636 21576
rect 27430 21564 27436 21576
rect 27488 21564 27494 21616
rect 30558 21604 30564 21616
rect 30519 21576 30564 21604
rect 30558 21564 30564 21576
rect 30616 21604 30622 21616
rect 31938 21604 31944 21616
rect 30616 21576 31944 21604
rect 30616 21564 30622 21576
rect 31938 21564 31944 21576
rect 31996 21564 32002 21616
rect 35434 21604 35440 21616
rect 35360 21576 35440 21604
rect 25593 21539 25651 21545
rect 25593 21536 25605 21539
rect 25096 21508 25605 21536
rect 25096 21496 25102 21508
rect 25593 21505 25605 21508
rect 25639 21505 25651 21539
rect 25593 21499 25651 21505
rect 26050 21496 26056 21548
rect 26108 21536 26114 21548
rect 26237 21539 26295 21545
rect 26237 21536 26249 21539
rect 26108 21508 26249 21536
rect 26108 21496 26114 21508
rect 26237 21505 26249 21508
rect 26283 21505 26295 21539
rect 26418 21536 26424 21548
rect 26379 21508 26424 21536
rect 26237 21499 26295 21505
rect 26418 21496 26424 21508
rect 26476 21496 26482 21548
rect 28074 21536 28080 21548
rect 28035 21508 28080 21536
rect 28074 21496 28080 21508
rect 28132 21496 28138 21548
rect 30006 21536 30012 21548
rect 29967 21508 30012 21536
rect 30006 21496 30012 21508
rect 30064 21496 30070 21548
rect 30466 21536 30472 21548
rect 30427 21508 30472 21536
rect 30466 21496 30472 21508
rect 30524 21496 30530 21548
rect 30650 21536 30656 21548
rect 30611 21508 30656 21536
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 31110 21496 31116 21548
rect 31168 21536 31174 21548
rect 31665 21539 31723 21545
rect 31665 21536 31677 21539
rect 31168 21508 31677 21536
rect 31168 21496 31174 21508
rect 31665 21505 31677 21508
rect 31711 21505 31723 21539
rect 31665 21499 31723 21505
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 22244 21440 22477 21468
rect 22244 21428 22250 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 23382 21468 23388 21480
rect 23343 21440 23388 21468
rect 22465 21431 22523 21437
rect 23382 21428 23388 21440
rect 23440 21428 23446 21480
rect 27706 21428 27712 21480
rect 27764 21468 27770 21480
rect 27985 21471 28043 21477
rect 27985 21468 27997 21471
rect 27764 21440 27997 21468
rect 27764 21428 27770 21440
rect 27985 21437 27997 21440
rect 28031 21437 28043 21471
rect 27985 21431 28043 21437
rect 31294 21428 31300 21480
rect 31352 21468 31358 21480
rect 31481 21471 31539 21477
rect 31481 21468 31493 21471
rect 31352 21440 31493 21468
rect 31352 21428 31358 21440
rect 31481 21437 31493 21440
rect 31527 21437 31539 21471
rect 31481 21431 31539 21437
rect 26053 21403 26111 21409
rect 26053 21369 26065 21403
rect 26099 21369 26111 21403
rect 31680 21400 31708 21499
rect 31754 21496 31760 21548
rect 31812 21536 31818 21548
rect 31812 21508 31905 21536
rect 31812 21496 31818 21508
rect 32214 21496 32220 21548
rect 32272 21536 32278 21548
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 32272 21508 32321 21536
rect 32272 21496 32278 21508
rect 32309 21505 32321 21508
rect 32355 21505 32367 21539
rect 33686 21536 33692 21548
rect 33647 21508 33692 21536
rect 32309 21499 32367 21505
rect 33686 21496 33692 21508
rect 33744 21496 33750 21548
rect 35360 21545 35388 21576
rect 35434 21564 35440 21576
rect 35492 21564 35498 21616
rect 35713 21607 35771 21613
rect 35713 21573 35725 21607
rect 35759 21604 35771 21607
rect 35759 21576 40540 21604
rect 35759 21573 35771 21576
rect 35713 21567 35771 21573
rect 33873 21539 33931 21545
rect 33873 21505 33885 21539
rect 33919 21505 33931 21539
rect 33873 21499 33931 21505
rect 35345 21539 35403 21545
rect 35345 21505 35357 21539
rect 35391 21505 35403 21539
rect 35526 21536 35532 21548
rect 35487 21508 35532 21536
rect 35345 21499 35403 21505
rect 31772 21468 31800 21496
rect 32582 21468 32588 21480
rect 31772 21440 32588 21468
rect 32582 21428 32588 21440
rect 32640 21428 32646 21480
rect 32950 21428 32956 21480
rect 33008 21468 33014 21480
rect 33137 21471 33195 21477
rect 33137 21468 33149 21471
rect 33008 21440 33149 21468
rect 33008 21428 33014 21440
rect 33137 21437 33149 21440
rect 33183 21468 33195 21471
rect 33888 21468 33916 21499
rect 35526 21496 35532 21508
rect 35584 21496 35590 21548
rect 35894 21496 35900 21548
rect 35952 21536 35958 21548
rect 36449 21539 36507 21545
rect 36449 21536 36461 21539
rect 35952 21508 36461 21536
rect 35952 21496 35958 21508
rect 36449 21505 36461 21508
rect 36495 21505 36507 21539
rect 36630 21536 36636 21548
rect 36591 21508 36636 21536
rect 36449 21499 36507 21505
rect 36630 21496 36636 21508
rect 36688 21496 36694 21548
rect 37366 21496 37372 21548
rect 37424 21536 37430 21548
rect 37645 21539 37703 21545
rect 37645 21536 37657 21539
rect 37424 21508 37657 21536
rect 37424 21496 37430 21508
rect 37645 21505 37657 21508
rect 37691 21505 37703 21539
rect 38194 21536 38200 21548
rect 37645 21499 37703 21505
rect 38028 21508 38200 21536
rect 34425 21471 34483 21477
rect 34425 21468 34437 21471
rect 33183 21440 34437 21468
rect 33183 21437 33195 21440
rect 33137 21431 33195 21437
rect 34425 21437 34437 21440
rect 34471 21468 34483 21471
rect 36648 21468 36676 21496
rect 37550 21468 37556 21480
rect 34471 21440 36676 21468
rect 37511 21440 37556 21468
rect 34471 21437 34483 21440
rect 34425 21431 34483 21437
rect 37550 21428 37556 21440
rect 37608 21428 37614 21480
rect 38028 21477 38056 21508
rect 38194 21496 38200 21508
rect 38252 21536 38258 21548
rect 40512 21545 40540 21576
rect 40678 21564 40684 21616
rect 40736 21604 40742 21616
rect 42058 21604 42064 21616
rect 40736 21576 42064 21604
rect 40736 21564 40742 21576
rect 42058 21564 42064 21576
rect 42116 21564 42122 21616
rect 42150 21564 42156 21616
rect 42208 21604 42214 21616
rect 43714 21604 43720 21616
rect 42208 21576 42840 21604
rect 43675 21576 43720 21604
rect 42208 21564 42214 21576
rect 38657 21539 38715 21545
rect 38657 21536 38669 21539
rect 38252 21508 38669 21536
rect 38252 21496 38258 21508
rect 38657 21505 38669 21508
rect 38703 21505 38715 21539
rect 38657 21499 38715 21505
rect 40497 21539 40555 21545
rect 40497 21505 40509 21539
rect 40543 21505 40555 21539
rect 40497 21499 40555 21505
rect 40586 21496 40592 21548
rect 40644 21536 40650 21548
rect 41141 21539 41199 21545
rect 41141 21536 41153 21539
rect 40644 21508 41153 21536
rect 40644 21496 40650 21508
rect 41141 21505 41153 21508
rect 41187 21505 41199 21539
rect 42705 21539 42763 21545
rect 42705 21536 42717 21539
rect 41141 21499 41199 21505
rect 41386 21508 42717 21536
rect 38013 21471 38071 21477
rect 38013 21437 38025 21471
rect 38059 21437 38071 21471
rect 38013 21431 38071 21437
rect 38470 21428 38476 21480
rect 38528 21468 38534 21480
rect 38565 21471 38623 21477
rect 38565 21468 38577 21471
rect 38528 21440 38577 21468
rect 38528 21428 38534 21440
rect 38565 21437 38577 21440
rect 38611 21437 38623 21471
rect 38565 21431 38623 21437
rect 41046 21428 41052 21480
rect 41104 21468 41110 21480
rect 41386 21468 41414 21508
rect 42705 21505 42717 21508
rect 42751 21505 42763 21539
rect 42812 21522 42840 21576
rect 43714 21564 43720 21576
rect 43772 21564 43778 21616
rect 44450 21564 44456 21616
rect 44508 21604 44514 21616
rect 44821 21607 44879 21613
rect 44821 21604 44833 21607
rect 44508 21576 44833 21604
rect 44508 21564 44514 21576
rect 44821 21573 44833 21576
rect 44867 21573 44879 21607
rect 44821 21567 44879 21573
rect 45278 21564 45284 21616
rect 45336 21564 45342 21616
rect 46566 21564 46572 21616
rect 46624 21604 46630 21616
rect 54478 21604 54484 21616
rect 46624 21576 54484 21604
rect 46624 21564 46630 21576
rect 47762 21536 47768 21548
rect 47723 21508 47768 21536
rect 42705 21499 42763 21505
rect 47762 21496 47768 21508
rect 47820 21496 47826 21548
rect 47854 21496 47860 21548
rect 47912 21536 47918 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47912 21508 47961 21536
rect 47912 21496 47918 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 48222 21496 48228 21548
rect 48280 21536 48286 21548
rect 48961 21539 49019 21545
rect 48961 21536 48973 21539
rect 48280 21508 48973 21536
rect 48280 21496 48286 21508
rect 48961 21505 48973 21508
rect 49007 21505 49019 21539
rect 48961 21499 49019 21505
rect 49234 21496 49240 21548
rect 49292 21536 49298 21548
rect 54128 21545 54156 21576
rect 54478 21564 54484 21576
rect 54536 21564 54542 21616
rect 49329 21539 49387 21545
rect 49329 21536 49341 21539
rect 49292 21508 49341 21536
rect 49292 21496 49298 21508
rect 49329 21505 49341 21508
rect 49375 21505 49387 21539
rect 49329 21499 49387 21505
rect 54113 21539 54171 21545
rect 54113 21505 54125 21539
rect 54159 21505 54171 21539
rect 54386 21536 54392 21548
rect 54347 21508 54392 21536
rect 54113 21499 54171 21505
rect 54386 21496 54392 21508
rect 54444 21496 54450 21548
rect 54573 21539 54631 21545
rect 54573 21505 54585 21539
rect 54619 21536 54631 21539
rect 55030 21536 55036 21548
rect 54619 21508 55036 21536
rect 54619 21505 54631 21508
rect 54573 21499 54631 21505
rect 55030 21496 55036 21508
rect 55088 21496 55094 21548
rect 55214 21536 55220 21548
rect 55175 21508 55220 21536
rect 55214 21496 55220 21508
rect 55272 21496 55278 21548
rect 56870 21536 56876 21548
rect 56831 21508 56876 21536
rect 56870 21496 56876 21508
rect 56928 21496 56934 21548
rect 56962 21496 56968 21548
rect 57020 21536 57026 21548
rect 57057 21539 57115 21545
rect 57057 21536 57069 21539
rect 57020 21508 57069 21536
rect 57020 21496 57026 21508
rect 57057 21505 57069 21508
rect 57103 21505 57115 21539
rect 57057 21499 57115 21505
rect 57882 21496 57888 21548
rect 57940 21536 57946 21548
rect 58069 21539 58127 21545
rect 58069 21536 58081 21539
rect 57940 21508 58081 21536
rect 57940 21496 57946 21508
rect 58069 21505 58081 21508
rect 58115 21505 58127 21539
rect 58069 21499 58127 21505
rect 58253 21539 58311 21545
rect 58253 21505 58265 21539
rect 58299 21536 58311 21539
rect 58342 21536 58348 21548
rect 58299 21508 58348 21536
rect 58299 21505 58311 21508
rect 58253 21499 58311 21505
rect 58342 21496 58348 21508
rect 58400 21496 58406 21548
rect 41104 21440 41414 21468
rect 41104 21428 41110 21440
rect 43438 21428 43444 21480
rect 43496 21468 43502 21480
rect 44545 21471 44603 21477
rect 44545 21468 44557 21471
rect 43496 21440 44557 21468
rect 43496 21428 43502 21440
rect 44545 21437 44557 21440
rect 44591 21468 44603 21471
rect 44591 21440 46980 21468
rect 44591 21437 44603 21440
rect 44545 21431 44603 21437
rect 32306 21400 32312 21412
rect 31680 21372 32312 21400
rect 26053 21363 26111 21369
rect 25498 21332 25504 21344
rect 25459 21304 25504 21332
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 25682 21292 25688 21344
rect 25740 21332 25746 21344
rect 26068 21332 26096 21363
rect 32306 21360 32312 21372
rect 32364 21400 32370 21412
rect 32401 21403 32459 21409
rect 32401 21400 32413 21403
rect 32364 21372 32413 21400
rect 32364 21360 32370 21372
rect 32401 21369 32413 21372
rect 32447 21369 32459 21403
rect 32401 21363 32459 21369
rect 46952 21344 46980 21440
rect 27249 21335 27307 21341
rect 27249 21332 27261 21335
rect 25740 21304 27261 21332
rect 25740 21292 25746 21304
rect 27249 21301 27261 21304
rect 27295 21332 27307 21335
rect 28626 21332 28632 21344
rect 27295 21304 28632 21332
rect 27295 21301 27307 21304
rect 27249 21295 27307 21301
rect 28626 21292 28632 21304
rect 28684 21332 28690 21344
rect 32950 21332 32956 21344
rect 28684 21304 32956 21332
rect 28684 21292 28690 21304
rect 32950 21292 32956 21304
rect 33008 21292 33014 21344
rect 33778 21332 33784 21344
rect 33739 21304 33784 21332
rect 33778 21292 33784 21304
rect 33836 21292 33842 21344
rect 43162 21292 43168 21344
rect 43220 21332 43226 21344
rect 46293 21335 46351 21341
rect 46293 21332 46305 21335
rect 43220 21304 46305 21332
rect 43220 21292 43226 21304
rect 46293 21301 46305 21304
rect 46339 21301 46351 21335
rect 46934 21332 46940 21344
rect 46895 21304 46940 21332
rect 46293 21295 46351 21301
rect 46934 21292 46940 21304
rect 46992 21292 46998 21344
rect 48958 21332 48964 21344
rect 48919 21304 48964 21332
rect 48958 21292 48964 21304
rect 49016 21292 49022 21344
rect 54205 21335 54263 21341
rect 54205 21301 54217 21335
rect 54251 21332 54263 21335
rect 54570 21332 54576 21344
rect 54251 21304 54576 21332
rect 54251 21301 54263 21304
rect 54205 21295 54263 21301
rect 54570 21292 54576 21304
rect 54628 21292 54634 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 23658 21128 23664 21140
rect 23619 21100 23664 21128
rect 23658 21088 23664 21100
rect 23716 21088 23722 21140
rect 24581 21131 24639 21137
rect 24581 21097 24593 21131
rect 24627 21128 24639 21131
rect 24670 21128 24676 21140
rect 24627 21100 24676 21128
rect 24627 21097 24639 21100
rect 24581 21091 24639 21097
rect 23842 20924 23848 20936
rect 23803 20896 23848 20924
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 24029 20927 24087 20933
rect 24029 20893 24041 20927
rect 24075 20924 24087 20927
rect 24596 20924 24624 21091
rect 24670 21088 24676 21100
rect 24728 21088 24734 21140
rect 24765 21131 24823 21137
rect 24765 21097 24777 21131
rect 24811 21128 24823 21131
rect 24946 21128 24952 21140
rect 24811 21100 24952 21128
rect 24811 21097 24823 21100
rect 24765 21091 24823 21097
rect 24946 21088 24952 21100
rect 25004 21128 25010 21140
rect 25961 21131 26019 21137
rect 25961 21128 25973 21131
rect 25004 21100 25973 21128
rect 25004 21088 25010 21100
rect 25961 21097 25973 21100
rect 26007 21097 26019 21131
rect 25961 21091 26019 21097
rect 27801 21131 27859 21137
rect 27801 21097 27813 21131
rect 27847 21128 27859 21131
rect 27890 21128 27896 21140
rect 27847 21100 27896 21128
rect 27847 21097 27859 21100
rect 27801 21091 27859 21097
rect 27890 21088 27896 21100
rect 27948 21088 27954 21140
rect 27985 21131 28043 21137
rect 27985 21097 27997 21131
rect 28031 21128 28043 21131
rect 28074 21128 28080 21140
rect 28031 21100 28080 21128
rect 28031 21097 28043 21100
rect 27985 21091 28043 21097
rect 28074 21088 28080 21100
rect 28132 21088 28138 21140
rect 29825 21131 29883 21137
rect 29825 21097 29837 21131
rect 29871 21128 29883 21131
rect 30282 21128 30288 21140
rect 29871 21100 30288 21128
rect 29871 21097 29883 21100
rect 29825 21091 29883 21097
rect 30282 21088 30288 21100
rect 30340 21088 30346 21140
rect 31478 21128 31484 21140
rect 31439 21100 31484 21128
rect 31478 21088 31484 21100
rect 31536 21088 31542 21140
rect 32306 21128 32312 21140
rect 32267 21100 32312 21128
rect 32306 21088 32312 21100
rect 32364 21088 32370 21140
rect 33137 21131 33195 21137
rect 33137 21097 33149 21131
rect 33183 21097 33195 21131
rect 33318 21128 33324 21140
rect 33279 21100 33324 21128
rect 33137 21091 33195 21097
rect 31665 21063 31723 21069
rect 31665 21060 31677 21063
rect 30668 21032 31677 21060
rect 30668 21004 30696 21032
rect 31665 21029 31677 21032
rect 31711 21029 31723 21063
rect 33152 21060 33180 21091
rect 33318 21088 33324 21100
rect 33376 21088 33382 21140
rect 35894 21128 35900 21140
rect 35855 21100 35900 21128
rect 35894 21088 35900 21100
rect 35952 21088 35958 21140
rect 37553 21131 37611 21137
rect 37553 21097 37565 21131
rect 37599 21128 37611 21131
rect 38102 21128 38108 21140
rect 37599 21100 38108 21128
rect 37599 21097 37611 21100
rect 37553 21091 37611 21097
rect 38102 21088 38108 21100
rect 38160 21088 38166 21140
rect 38286 21088 38292 21140
rect 38344 21128 38350 21140
rect 38565 21131 38623 21137
rect 38565 21128 38577 21131
rect 38344 21100 38577 21128
rect 38344 21088 38350 21100
rect 38565 21097 38577 21100
rect 38611 21097 38623 21131
rect 38565 21091 38623 21097
rect 44637 21131 44695 21137
rect 44637 21097 44649 21131
rect 44683 21128 44695 21131
rect 45738 21128 45744 21140
rect 44683 21100 45744 21128
rect 44683 21097 44695 21100
rect 44637 21091 44695 21097
rect 45738 21088 45744 21100
rect 45796 21088 45802 21140
rect 45833 21131 45891 21137
rect 45833 21097 45845 21131
rect 45879 21128 45891 21131
rect 46934 21128 46940 21140
rect 45879 21100 46940 21128
rect 45879 21097 45891 21100
rect 45833 21091 45891 21097
rect 46934 21088 46940 21100
rect 46992 21088 46998 21140
rect 48869 21131 48927 21137
rect 48869 21097 48881 21131
rect 48915 21128 48927 21131
rect 49142 21128 49148 21140
rect 48915 21100 49148 21128
rect 48915 21097 48927 21100
rect 48869 21091 48927 21097
rect 49142 21088 49148 21100
rect 49200 21088 49206 21140
rect 54113 21131 54171 21137
rect 54113 21097 54125 21131
rect 54159 21128 54171 21131
rect 54386 21128 54392 21140
rect 54159 21100 54392 21128
rect 54159 21097 54171 21100
rect 54113 21091 54171 21097
rect 54386 21088 54392 21100
rect 54444 21088 54450 21140
rect 56870 21128 56876 21140
rect 56831 21100 56876 21128
rect 56870 21088 56876 21100
rect 56928 21088 56934 21140
rect 56962 21088 56968 21140
rect 57020 21128 57026 21140
rect 57701 21131 57759 21137
rect 57701 21128 57713 21131
rect 57020 21100 57713 21128
rect 57020 21088 57026 21100
rect 57701 21097 57713 21100
rect 57747 21097 57759 21131
rect 57882 21128 57888 21140
rect 57843 21100 57888 21128
rect 57701 21091 57759 21097
rect 57882 21088 57888 21100
rect 57940 21088 57946 21140
rect 33686 21060 33692 21072
rect 33152 21032 33692 21060
rect 31665 21023 31723 21029
rect 26050 20952 26056 21004
rect 26108 20992 26114 21004
rect 26237 20995 26295 21001
rect 26237 20992 26249 20995
rect 26108 20964 26249 20992
rect 26108 20952 26114 20964
rect 26237 20961 26249 20964
rect 26283 20961 26295 20995
rect 26237 20955 26295 20961
rect 27706 20952 27712 21004
rect 27764 20992 27770 21004
rect 28537 20995 28595 21001
rect 28537 20992 28549 20995
rect 27764 20964 28549 20992
rect 27764 20952 27770 20964
rect 28537 20961 28549 20964
rect 28583 20961 28595 20995
rect 28721 20995 28779 21001
rect 28721 20992 28733 20995
rect 28537 20955 28595 20961
rect 28644 20964 28733 20992
rect 26142 20924 26148 20936
rect 24075 20896 24624 20924
rect 26103 20896 26148 20924
rect 24075 20893 24087 20896
rect 24029 20887 24087 20893
rect 26142 20884 26148 20896
rect 26200 20884 26206 20936
rect 26329 20927 26387 20933
rect 26329 20893 26341 20927
rect 26375 20893 26387 20927
rect 26329 20887 26387 20893
rect 24762 20865 24768 20868
rect 24749 20859 24768 20865
rect 24749 20825 24761 20859
rect 24749 20819 24768 20825
rect 24762 20816 24768 20819
rect 24820 20816 24826 20868
rect 24854 20816 24860 20868
rect 24912 20856 24918 20868
rect 24949 20859 25007 20865
rect 24949 20856 24961 20859
rect 24912 20828 24961 20856
rect 24912 20816 24918 20828
rect 24949 20825 24961 20828
rect 24995 20825 25007 20859
rect 24949 20819 25007 20825
rect 25498 20816 25504 20868
rect 25556 20856 25562 20868
rect 26344 20856 26372 20887
rect 26418 20884 26424 20936
rect 26476 20924 26482 20936
rect 28442 20924 28448 20936
rect 26476 20896 27752 20924
rect 28403 20896 28448 20924
rect 26476 20884 26482 20896
rect 27617 20859 27675 20865
rect 27617 20856 27629 20859
rect 25556 20828 27629 20856
rect 25556 20816 25562 20828
rect 27617 20825 27629 20828
rect 27663 20825 27675 20859
rect 27724 20856 27752 20896
rect 28442 20884 28448 20896
rect 28500 20884 28506 20936
rect 28534 20856 28540 20868
rect 27724 20828 28540 20856
rect 27617 20819 27675 20825
rect 28534 20816 28540 20828
rect 28592 20816 28598 20868
rect 27798 20748 27804 20800
rect 27856 20797 27862 20800
rect 27856 20791 27875 20797
rect 27863 20788 27875 20791
rect 28644 20788 28672 20964
rect 28721 20961 28733 20964
rect 28767 20961 28779 20995
rect 30650 20992 30656 21004
rect 28721 20955 28779 20961
rect 30208 20964 30656 20992
rect 30006 20924 30012 20936
rect 29919 20896 30012 20924
rect 30006 20884 30012 20896
rect 30064 20884 30070 20936
rect 30208 20933 30236 20964
rect 30650 20952 30656 20964
rect 30708 20952 30714 21004
rect 30926 20952 30932 21004
rect 30984 20992 30990 21004
rect 30984 20964 31524 20992
rect 30984 20952 30990 20964
rect 30193 20927 30251 20933
rect 30193 20893 30205 20927
rect 30239 20893 30251 20927
rect 30193 20887 30251 20893
rect 30285 20927 30343 20933
rect 30285 20893 30297 20927
rect 30331 20924 30343 20927
rect 30466 20924 30472 20936
rect 30331 20896 30472 20924
rect 30331 20893 30343 20896
rect 30285 20887 30343 20893
rect 30466 20884 30472 20896
rect 30524 20884 30530 20936
rect 31294 20884 31300 20936
rect 31352 20924 31358 20936
rect 31496 20933 31524 20964
rect 31389 20927 31447 20933
rect 31389 20924 31401 20927
rect 31352 20896 31401 20924
rect 31352 20884 31358 20896
rect 31389 20893 31401 20896
rect 31435 20893 31447 20927
rect 31389 20887 31447 20893
rect 31481 20927 31539 20933
rect 31481 20893 31493 20927
rect 31527 20924 31539 20927
rect 31570 20924 31576 20936
rect 31527 20896 31576 20924
rect 31527 20893 31539 20896
rect 31481 20887 31539 20893
rect 28721 20859 28779 20865
rect 28721 20825 28733 20859
rect 28767 20856 28779 20859
rect 30024 20856 30052 20884
rect 28767 20828 30052 20856
rect 28767 20825 28779 20828
rect 28721 20819 28779 20825
rect 30558 20816 30564 20868
rect 30616 20856 30622 20868
rect 31205 20859 31263 20865
rect 31205 20856 31217 20859
rect 30616 20828 31217 20856
rect 30616 20816 30622 20828
rect 31205 20825 31217 20828
rect 31251 20825 31263 20859
rect 31205 20819 31263 20825
rect 27863 20760 28672 20788
rect 31404 20788 31432 20887
rect 31570 20884 31576 20896
rect 31628 20884 31634 20936
rect 31680 20924 31708 21023
rect 33686 21020 33692 21032
rect 33744 21020 33750 21072
rect 34149 21063 34207 21069
rect 34149 21029 34161 21063
rect 34195 21060 34207 21063
rect 35526 21060 35532 21072
rect 34195 21032 35532 21060
rect 34195 21029 34207 21032
rect 34149 21023 34207 21029
rect 35526 21020 35532 21032
rect 35584 21020 35590 21072
rect 41509 21063 41567 21069
rect 41509 21029 41521 21063
rect 41555 21060 41567 21063
rect 42337 21063 42395 21069
rect 42337 21060 42349 21063
rect 41555 21032 42349 21060
rect 41555 21029 41567 21032
rect 41509 21023 41567 21029
rect 42337 21029 42349 21032
rect 42383 21060 42395 21063
rect 42426 21060 42432 21072
rect 42383 21032 42432 21060
rect 42383 21029 42395 21032
rect 42337 21023 42395 21029
rect 42426 21020 42432 21032
rect 42484 21020 42490 21072
rect 47486 21060 47492 21072
rect 47447 21032 47492 21060
rect 47486 21020 47492 21032
rect 47544 21020 47550 21072
rect 52546 21060 52552 21072
rect 52507 21032 52552 21060
rect 52546 21020 52552 21032
rect 52604 21020 52610 21072
rect 55490 21060 55496 21072
rect 53392 21032 55496 21060
rect 33778 20952 33784 21004
rect 33836 20992 33842 21004
rect 33965 20995 34023 21001
rect 33965 20992 33977 20995
rect 33836 20964 33977 20992
rect 33836 20952 33842 20964
rect 33965 20961 33977 20964
rect 34011 20961 34023 20995
rect 33965 20955 34023 20961
rect 35621 20995 35679 21001
rect 35621 20961 35633 20995
rect 35667 20992 35679 20995
rect 35710 20992 35716 21004
rect 35667 20964 35716 20992
rect 35667 20961 35679 20964
rect 35621 20955 35679 20961
rect 35710 20952 35716 20964
rect 35768 20952 35774 21004
rect 38194 20992 38200 21004
rect 38155 20964 38200 20992
rect 38194 20952 38200 20964
rect 38252 20952 38258 21004
rect 41969 20995 42027 21001
rect 41969 20961 41981 20995
rect 42015 20992 42027 20995
rect 42889 20995 42947 21001
rect 42889 20992 42901 20995
rect 42015 20964 42901 20992
rect 42015 20961 42027 20964
rect 41969 20955 42027 20961
rect 42889 20961 42901 20964
rect 42935 20992 42947 20995
rect 43254 20992 43260 21004
rect 42935 20964 43260 20992
rect 42935 20961 42947 20964
rect 42889 20955 42947 20961
rect 43254 20952 43260 20964
rect 43312 20952 43318 21004
rect 47213 20995 47271 21001
rect 47213 20961 47225 20995
rect 47259 20992 47271 20995
rect 48041 20995 48099 21001
rect 48041 20992 48053 20995
rect 47259 20964 48053 20992
rect 47259 20961 47271 20964
rect 47213 20955 47271 20961
rect 48041 20961 48053 20964
rect 48087 20961 48099 20995
rect 48041 20955 48099 20961
rect 51258 20952 51264 21004
rect 51316 20992 51322 21004
rect 51994 20992 52000 21004
rect 51316 20964 52000 20992
rect 51316 20952 51322 20964
rect 51994 20952 52000 20964
rect 52052 20992 52058 21004
rect 52089 20995 52147 21001
rect 52089 20992 52101 20995
rect 52052 20964 52101 20992
rect 52052 20952 52058 20964
rect 52089 20961 52101 20964
rect 52135 20961 52147 20995
rect 52564 20992 52592 21020
rect 52564 20964 53144 20992
rect 52089 20955 52147 20961
rect 32217 20927 32275 20933
rect 32217 20924 32229 20927
rect 31680 20896 32229 20924
rect 32217 20893 32229 20896
rect 32263 20893 32275 20927
rect 32217 20887 32275 20893
rect 34149 20927 34207 20933
rect 34149 20893 34161 20927
rect 34195 20924 34207 20927
rect 34514 20924 34520 20936
rect 34195 20896 34520 20924
rect 34195 20893 34207 20896
rect 34149 20887 34207 20893
rect 34514 20884 34520 20896
rect 34572 20884 34578 20936
rect 35526 20924 35532 20936
rect 35487 20896 35532 20924
rect 35526 20884 35532 20896
rect 35584 20884 35590 20936
rect 37366 20924 37372 20936
rect 35636 20896 37372 20924
rect 32950 20856 32956 20868
rect 32911 20828 32956 20856
rect 32950 20816 32956 20828
rect 33008 20816 33014 20868
rect 33169 20859 33227 20865
rect 33169 20825 33181 20859
rect 33215 20856 33227 20859
rect 33502 20856 33508 20868
rect 33215 20828 33508 20856
rect 33215 20825 33227 20828
rect 33169 20819 33227 20825
rect 33502 20816 33508 20828
rect 33560 20856 33566 20868
rect 33781 20859 33839 20865
rect 33781 20856 33793 20859
rect 33560 20828 33793 20856
rect 33560 20816 33566 20828
rect 33781 20825 33793 20828
rect 33827 20825 33839 20859
rect 33781 20819 33839 20825
rect 35636 20800 35664 20896
rect 37366 20884 37372 20896
rect 37424 20884 37430 20936
rect 37550 20924 37556 20936
rect 37511 20896 37556 20924
rect 37550 20884 37556 20896
rect 37608 20884 37614 20936
rect 38381 20927 38439 20933
rect 38381 20893 38393 20927
rect 38427 20924 38439 20927
rect 38470 20924 38476 20936
rect 38427 20896 38476 20924
rect 38427 20893 38439 20896
rect 38381 20887 38439 20893
rect 38470 20884 38476 20896
rect 38528 20884 38534 20936
rect 42426 20884 42432 20936
rect 42484 20884 42490 20936
rect 47121 20927 47179 20933
rect 47121 20893 47133 20927
rect 47167 20893 47179 20927
rect 47946 20924 47952 20936
rect 47907 20896 47952 20924
rect 47121 20887 47179 20893
rect 42444 20856 42472 20884
rect 43162 20856 43168 20868
rect 42444 20828 43024 20856
rect 43123 20828 43168 20856
rect 32214 20788 32220 20800
rect 31404 20760 32220 20788
rect 27863 20757 27875 20760
rect 27856 20751 27875 20757
rect 27856 20748 27862 20751
rect 32214 20748 32220 20760
rect 32272 20748 32278 20800
rect 35618 20748 35624 20800
rect 35676 20748 35682 20800
rect 36449 20791 36507 20797
rect 36449 20757 36461 20791
rect 36495 20788 36507 20791
rect 36630 20788 36636 20800
rect 36495 20760 36636 20788
rect 36495 20757 36507 20760
rect 36449 20751 36507 20757
rect 36630 20748 36636 20760
rect 36688 20788 36694 20800
rect 39390 20788 39396 20800
rect 36688 20760 39396 20788
rect 36688 20748 36694 20760
rect 39390 20748 39396 20760
rect 39448 20748 39454 20800
rect 42429 20791 42487 20797
rect 42429 20757 42441 20791
rect 42475 20788 42487 20791
rect 42610 20788 42616 20800
rect 42475 20760 42616 20788
rect 42475 20757 42487 20760
rect 42429 20751 42487 20757
rect 42610 20748 42616 20760
rect 42668 20748 42674 20800
rect 42996 20788 43024 20828
rect 43162 20816 43168 20828
rect 43220 20816 43226 20868
rect 47136 20856 47164 20887
rect 47946 20884 47952 20896
rect 48004 20884 48010 20936
rect 48130 20924 48136 20936
rect 48091 20896 48136 20924
rect 48130 20884 48136 20896
rect 48188 20884 48194 20936
rect 48222 20884 48228 20936
rect 48280 20924 48286 20936
rect 48685 20927 48743 20933
rect 48685 20924 48697 20927
rect 48280 20896 48697 20924
rect 48280 20884 48286 20896
rect 48685 20893 48697 20896
rect 48731 20893 48743 20927
rect 48685 20887 48743 20893
rect 48869 20927 48927 20933
rect 48869 20893 48881 20927
rect 48915 20924 48927 20927
rect 48958 20924 48964 20936
rect 48915 20896 48964 20924
rect 48915 20893 48927 20896
rect 48869 20887 48927 20893
rect 48958 20884 48964 20896
rect 49016 20884 49022 20936
rect 49142 20924 49148 20936
rect 49103 20896 49148 20924
rect 49142 20884 49148 20896
rect 49200 20884 49206 20936
rect 50890 20884 50896 20936
rect 50948 20924 50954 20936
rect 50985 20927 51043 20933
rect 50985 20924 50997 20927
rect 50948 20896 50997 20924
rect 50948 20884 50954 20896
rect 50985 20893 50997 20896
rect 51031 20893 51043 20927
rect 51350 20924 51356 20936
rect 51311 20896 51356 20924
rect 50985 20887 51043 20893
rect 51350 20884 51356 20896
rect 51408 20884 51414 20936
rect 51534 20884 51540 20936
rect 51592 20924 51598 20936
rect 52181 20927 52239 20933
rect 52181 20924 52193 20927
rect 51592 20896 52193 20924
rect 51592 20884 51598 20896
rect 52181 20893 52193 20896
rect 52227 20893 52239 20927
rect 53006 20924 53012 20936
rect 52967 20896 53012 20924
rect 52181 20887 52239 20893
rect 53006 20884 53012 20896
rect 53064 20884 53070 20936
rect 53116 20933 53144 20964
rect 53101 20927 53159 20933
rect 53101 20893 53113 20927
rect 53147 20893 53159 20927
rect 53282 20924 53288 20936
rect 53243 20896 53288 20924
rect 53101 20887 53159 20893
rect 53282 20884 53288 20896
rect 53340 20884 53346 20936
rect 47394 20856 47400 20868
rect 43364 20828 43654 20856
rect 47136 20828 47400 20856
rect 43364 20788 43392 20828
rect 47394 20816 47400 20828
rect 47452 20856 47458 20868
rect 48240 20856 48268 20884
rect 47452 20828 48268 20856
rect 47452 20816 47458 20828
rect 44542 20788 44548 20800
rect 42996 20760 44548 20788
rect 44542 20748 44548 20760
rect 44600 20788 44606 20800
rect 45189 20791 45247 20797
rect 45189 20788 45201 20791
rect 44600 20760 45201 20788
rect 44600 20748 44606 20760
rect 45189 20757 45201 20760
rect 45235 20788 45247 20791
rect 45278 20788 45284 20800
rect 45235 20760 45284 20788
rect 45235 20757 45247 20760
rect 45189 20751 45247 20757
rect 45278 20748 45284 20760
rect 45336 20748 45342 20800
rect 45738 20748 45744 20800
rect 45796 20788 45802 20800
rect 46293 20791 46351 20797
rect 46293 20788 46305 20791
rect 45796 20760 46305 20788
rect 45796 20748 45802 20760
rect 46293 20757 46305 20760
rect 46339 20757 46351 20791
rect 46293 20751 46351 20757
rect 51077 20791 51135 20797
rect 51077 20757 51089 20791
rect 51123 20788 51135 20791
rect 53392 20788 53420 21032
rect 55490 21020 55496 21032
rect 55548 21020 55554 21072
rect 55398 20952 55404 21004
rect 55456 20992 55462 21004
rect 55585 20995 55643 21001
rect 55585 20992 55597 20995
rect 55456 20964 55597 20992
rect 55456 20952 55462 20964
rect 55585 20961 55597 20964
rect 55631 20961 55643 20995
rect 55585 20955 55643 20961
rect 53834 20884 53840 20936
rect 53892 20924 53898 20936
rect 53929 20927 53987 20933
rect 53929 20924 53941 20927
rect 53892 20896 53941 20924
rect 53892 20884 53898 20896
rect 53929 20893 53941 20896
rect 53975 20924 53987 20927
rect 54018 20924 54024 20936
rect 53975 20896 54024 20924
rect 53975 20893 53987 20896
rect 53929 20887 53987 20893
rect 54018 20884 54024 20896
rect 54076 20884 54082 20936
rect 54294 20924 54300 20936
rect 54255 20896 54300 20924
rect 54294 20884 54300 20896
rect 54352 20884 54358 20936
rect 54389 20927 54447 20933
rect 54389 20893 54401 20927
rect 54435 20924 54447 20927
rect 54570 20924 54576 20936
rect 54435 20896 54576 20924
rect 54435 20893 54447 20896
rect 54389 20887 54447 20893
rect 54570 20884 54576 20896
rect 54628 20884 54634 20936
rect 55674 20924 55680 20936
rect 54956 20896 55680 20924
rect 53469 20859 53527 20865
rect 53469 20825 53481 20859
rect 53515 20856 53527 20859
rect 54956 20856 54984 20896
rect 55674 20884 55680 20896
rect 55732 20933 55738 20936
rect 55732 20927 55781 20933
rect 55732 20893 55735 20927
rect 55769 20893 55781 20927
rect 55732 20887 55781 20893
rect 55732 20884 55738 20887
rect 56502 20856 56508 20868
rect 53515 20828 54984 20856
rect 56463 20828 56508 20856
rect 53515 20825 53527 20828
rect 53469 20819 53527 20825
rect 56502 20816 56508 20828
rect 56560 20816 56566 20868
rect 56689 20859 56747 20865
rect 56689 20825 56701 20859
rect 56735 20825 56747 20859
rect 57514 20856 57520 20868
rect 57475 20828 57520 20856
rect 56689 20819 56747 20825
rect 51123 20760 53420 20788
rect 56045 20791 56103 20797
rect 51123 20757 51135 20760
rect 51077 20751 51135 20757
rect 56045 20757 56057 20791
rect 56091 20788 56103 20791
rect 56594 20788 56600 20800
rect 56091 20760 56600 20788
rect 56091 20757 56103 20760
rect 56045 20751 56103 20757
rect 56594 20748 56600 20760
rect 56652 20788 56658 20800
rect 56704 20788 56732 20819
rect 57514 20816 57520 20828
rect 57572 20816 57578 20868
rect 56652 20760 56732 20788
rect 56652 20748 56658 20760
rect 57698 20748 57704 20800
rect 57756 20797 57762 20800
rect 57756 20791 57775 20797
rect 57763 20757 57775 20791
rect 57756 20751 57775 20757
rect 57756 20748 57762 20751
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 24305 20587 24363 20593
rect 24305 20553 24317 20587
rect 24351 20584 24363 20587
rect 24762 20584 24768 20596
rect 24351 20556 24768 20584
rect 24351 20553 24363 20556
rect 24305 20547 24363 20553
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 25682 20584 25688 20596
rect 25643 20556 25688 20584
rect 25682 20544 25688 20556
rect 25740 20544 25746 20596
rect 26234 20584 26240 20596
rect 26195 20556 26240 20584
rect 26234 20544 26240 20556
rect 26292 20544 26298 20596
rect 26326 20544 26332 20596
rect 26384 20584 26390 20596
rect 26421 20587 26479 20593
rect 26421 20584 26433 20587
rect 26384 20556 26433 20584
rect 26384 20544 26390 20556
rect 26421 20553 26433 20556
rect 26467 20553 26479 20587
rect 26421 20547 26479 20553
rect 28077 20587 28135 20593
rect 28077 20553 28089 20587
rect 28123 20584 28135 20587
rect 28442 20584 28448 20596
rect 28123 20556 28448 20584
rect 28123 20553 28135 20556
rect 28077 20547 28135 20553
rect 28442 20544 28448 20556
rect 28500 20544 28506 20596
rect 28534 20544 28540 20596
rect 28592 20584 28598 20596
rect 29089 20587 29147 20593
rect 29089 20584 29101 20587
rect 28592 20556 29101 20584
rect 28592 20544 28598 20556
rect 29089 20553 29101 20556
rect 29135 20553 29147 20587
rect 30466 20584 30472 20596
rect 30427 20556 30472 20584
rect 29089 20547 29147 20553
rect 30466 20544 30472 20556
rect 30524 20544 30530 20596
rect 31478 20584 31484 20596
rect 31439 20556 31484 20584
rect 31478 20544 31484 20556
rect 31536 20544 31542 20596
rect 32493 20587 32551 20593
rect 32493 20584 32505 20587
rect 31588 20556 32505 20584
rect 22830 20516 22836 20528
rect 22791 20488 22836 20516
rect 22830 20476 22836 20488
rect 22888 20476 22894 20528
rect 23290 20476 23296 20528
rect 23348 20516 23354 20528
rect 25700 20516 25728 20544
rect 28626 20516 28632 20528
rect 23348 20488 25728 20516
rect 28587 20488 28632 20516
rect 23348 20476 23354 20488
rect 28626 20476 28632 20488
rect 28684 20476 28690 20528
rect 31294 20516 31300 20528
rect 30668 20488 31300 20516
rect 23492 20380 23520 20434
rect 23566 20408 23572 20460
rect 23624 20448 23630 20460
rect 23624 20420 23669 20448
rect 23624 20408 23630 20420
rect 24026 20408 24032 20460
rect 24084 20448 24090 20460
rect 24581 20451 24639 20457
rect 24581 20448 24593 20451
rect 24084 20420 24593 20448
rect 24084 20408 24090 20420
rect 24581 20417 24593 20420
rect 24627 20417 24639 20451
rect 24581 20411 24639 20417
rect 24673 20451 24731 20457
rect 24673 20417 24685 20451
rect 24719 20448 24731 20451
rect 25498 20448 25504 20460
rect 24719 20420 25504 20448
rect 24719 20417 24731 20420
rect 24673 20411 24731 20417
rect 25498 20408 25504 20420
rect 25556 20408 25562 20460
rect 26418 20408 26424 20460
rect 26476 20448 26482 20460
rect 26513 20451 26571 20457
rect 26513 20448 26525 20451
rect 26476 20420 26525 20448
rect 26476 20408 26482 20420
rect 26513 20417 26525 20420
rect 26559 20417 26571 20451
rect 26513 20411 26571 20417
rect 26602 20408 26608 20460
rect 26660 20448 26666 20460
rect 27890 20448 27896 20460
rect 26660 20420 26705 20448
rect 27851 20420 27896 20448
rect 26660 20408 26666 20420
rect 27890 20408 27896 20420
rect 27948 20408 27954 20460
rect 28077 20451 28135 20457
rect 28077 20417 28089 20451
rect 28123 20448 28135 20451
rect 28644 20448 28672 20476
rect 28123 20420 28672 20448
rect 29457 20451 29515 20457
rect 28123 20417 28135 20420
rect 28077 20411 28135 20417
rect 29457 20417 29469 20451
rect 29503 20448 29515 20451
rect 29730 20448 29736 20460
rect 29503 20420 29736 20448
rect 29503 20417 29515 20420
rect 29457 20411 29515 20417
rect 29730 20408 29736 20420
rect 29788 20408 29794 20460
rect 30469 20451 30527 20457
rect 30469 20417 30481 20451
rect 30515 20448 30527 20451
rect 30558 20448 30564 20460
rect 30515 20420 30564 20448
rect 30515 20417 30527 20420
rect 30469 20411 30527 20417
rect 30558 20408 30564 20420
rect 30616 20408 30622 20460
rect 30668 20457 30696 20488
rect 31294 20476 31300 20488
rect 31352 20476 31358 20528
rect 31588 20516 31616 20556
rect 32493 20553 32505 20556
rect 32539 20553 32551 20587
rect 32493 20547 32551 20553
rect 33686 20544 33692 20596
rect 33744 20584 33750 20596
rect 33781 20587 33839 20593
rect 33781 20584 33793 20587
rect 33744 20556 33793 20584
rect 33744 20544 33750 20556
rect 33781 20553 33793 20556
rect 33827 20553 33839 20587
rect 33781 20547 33839 20553
rect 34514 20544 34520 20596
rect 34572 20584 34578 20596
rect 35069 20587 35127 20593
rect 35069 20584 35081 20587
rect 34572 20556 35081 20584
rect 34572 20544 34578 20556
rect 35069 20553 35081 20556
rect 35115 20553 35127 20587
rect 35069 20547 35127 20553
rect 39209 20587 39267 20593
rect 39209 20553 39221 20587
rect 39255 20553 39267 20587
rect 41046 20584 41052 20596
rect 41007 20556 41052 20584
rect 39209 20547 39267 20553
rect 32677 20519 32735 20525
rect 32677 20516 32689 20519
rect 31404 20488 31616 20516
rect 31680 20488 32689 20516
rect 31404 20460 31432 20488
rect 31680 20460 31708 20488
rect 32677 20485 32689 20488
rect 32723 20485 32735 20519
rect 32677 20479 32735 20485
rect 30653 20451 30711 20457
rect 30653 20417 30665 20451
rect 30699 20417 30711 20451
rect 30926 20448 30932 20460
rect 30887 20420 30932 20448
rect 30653 20411 30711 20417
rect 30926 20408 30932 20420
rect 30984 20408 30990 20460
rect 31386 20448 31392 20460
rect 31347 20420 31392 20448
rect 31386 20408 31392 20420
rect 31444 20408 31450 20460
rect 31662 20448 31668 20460
rect 31623 20420 31668 20448
rect 31662 20408 31668 20420
rect 31720 20408 31726 20460
rect 31754 20408 31760 20460
rect 31812 20448 31818 20460
rect 32585 20451 32643 20457
rect 32585 20448 32597 20451
rect 31812 20420 32597 20448
rect 31812 20408 31818 20420
rect 32585 20417 32597 20420
rect 32631 20417 32643 20451
rect 32585 20411 32643 20417
rect 33226 20408 33232 20460
rect 33284 20448 33290 20460
rect 33321 20451 33379 20457
rect 33321 20448 33333 20451
rect 33284 20420 33333 20448
rect 33284 20408 33290 20420
rect 33321 20417 33333 20420
rect 33367 20417 33379 20451
rect 33321 20411 33379 20417
rect 33410 20408 33416 20460
rect 33468 20448 33474 20460
rect 33597 20451 33655 20457
rect 33468 20420 33513 20448
rect 33468 20408 33474 20420
rect 33597 20417 33609 20451
rect 33643 20448 33655 20451
rect 33778 20448 33784 20460
rect 33643 20420 33784 20448
rect 33643 20417 33655 20420
rect 33597 20411 33655 20417
rect 33778 20408 33784 20420
rect 33836 20408 33842 20460
rect 35434 20448 35440 20460
rect 35395 20420 35440 20448
rect 35434 20408 35440 20420
rect 35492 20408 35498 20460
rect 36633 20451 36691 20457
rect 36633 20417 36645 20451
rect 36679 20448 36691 20451
rect 36722 20448 36728 20460
rect 36679 20420 36728 20448
rect 36679 20417 36691 20420
rect 36633 20411 36691 20417
rect 36722 20408 36728 20420
rect 36780 20408 36786 20460
rect 36817 20451 36875 20457
rect 36817 20417 36829 20451
rect 36863 20448 36875 20451
rect 36906 20448 36912 20460
rect 36863 20420 36912 20448
rect 36863 20417 36875 20420
rect 36817 20411 36875 20417
rect 36906 20408 36912 20420
rect 36964 20408 36970 20460
rect 38838 20448 38844 20460
rect 38799 20420 38844 20448
rect 38838 20408 38844 20420
rect 38896 20408 38902 20460
rect 39224 20448 39252 20547
rect 41046 20544 41052 20556
rect 41104 20544 41110 20596
rect 43349 20587 43407 20593
rect 43349 20553 43361 20587
rect 43395 20584 43407 20587
rect 43438 20584 43444 20596
rect 43395 20556 43444 20584
rect 43395 20553 43407 20556
rect 43349 20547 43407 20553
rect 43438 20544 43444 20556
rect 43496 20544 43502 20596
rect 48409 20587 48467 20593
rect 48409 20553 48421 20587
rect 48455 20584 48467 20587
rect 48958 20584 48964 20596
rect 48455 20556 48964 20584
rect 48455 20553 48467 20556
rect 48409 20547 48467 20553
rect 48958 20544 48964 20556
rect 49016 20544 49022 20596
rect 53193 20587 53251 20593
rect 49252 20556 51074 20584
rect 46753 20519 46811 20525
rect 46753 20485 46765 20519
rect 46799 20516 46811 20519
rect 47946 20516 47952 20528
rect 46799 20488 47952 20516
rect 46799 20485 46811 20488
rect 46753 20479 46811 20485
rect 47946 20476 47952 20488
rect 48004 20516 48010 20528
rect 49252 20516 49280 20556
rect 51046 20528 51074 20556
rect 53193 20553 53205 20587
rect 53239 20584 53251 20587
rect 53282 20584 53288 20596
rect 53239 20556 53288 20584
rect 53239 20553 53251 20556
rect 53193 20547 53251 20553
rect 53282 20544 53288 20556
rect 53340 20544 53346 20596
rect 55214 20584 55220 20596
rect 54588 20556 55220 20584
rect 48004 20488 49280 20516
rect 48004 20476 48010 20488
rect 40034 20448 40040 20460
rect 39224 20420 40040 20448
rect 40034 20408 40040 20420
rect 40092 20448 40098 20460
rect 40221 20451 40279 20457
rect 40221 20448 40233 20451
rect 40092 20420 40233 20448
rect 40092 20408 40098 20420
rect 40221 20417 40233 20420
rect 40267 20417 40279 20451
rect 40221 20411 40279 20417
rect 41230 20408 41236 20460
rect 41288 20448 41294 20460
rect 41509 20451 41567 20457
rect 41509 20448 41521 20451
rect 41288 20420 41521 20448
rect 41288 20408 41294 20420
rect 41509 20417 41521 20420
rect 41555 20417 41567 20451
rect 41509 20411 41567 20417
rect 41690 20408 41696 20460
rect 41748 20448 41754 20460
rect 41874 20448 41880 20460
rect 41748 20420 41880 20448
rect 41748 20408 41754 20420
rect 41874 20408 41880 20420
rect 41932 20408 41938 20460
rect 42610 20448 42616 20460
rect 42571 20420 42616 20448
rect 42610 20408 42616 20420
rect 42668 20408 42674 20460
rect 44450 20448 44456 20460
rect 44411 20420 44456 20448
rect 44450 20408 44456 20420
rect 44508 20408 44514 20460
rect 45554 20448 45560 20460
rect 44836 20420 45560 20448
rect 24486 20380 24492 20392
rect 23492 20352 24492 20380
rect 24486 20340 24492 20352
rect 24544 20340 24550 20392
rect 24765 20383 24823 20389
rect 24765 20349 24777 20383
rect 24811 20349 24823 20383
rect 24765 20343 24823 20349
rect 26237 20383 26295 20389
rect 26237 20349 26249 20383
rect 26283 20349 26295 20383
rect 26237 20343 26295 20349
rect 23934 20272 23940 20324
rect 23992 20312 23998 20324
rect 24780 20312 24808 20343
rect 23992 20284 24808 20312
rect 26252 20312 26280 20343
rect 29270 20340 29276 20392
rect 29328 20380 29334 20392
rect 29365 20383 29423 20389
rect 29365 20380 29377 20383
rect 29328 20352 29377 20380
rect 29328 20340 29334 20352
rect 29365 20349 29377 20352
rect 29411 20349 29423 20383
rect 29365 20343 29423 20349
rect 30791 20383 30849 20389
rect 30791 20349 30803 20383
rect 30837 20380 30849 20383
rect 31478 20380 31484 20392
rect 30837 20352 31484 20380
rect 30837 20349 30849 20352
rect 30791 20343 30849 20349
rect 31478 20340 31484 20352
rect 31536 20340 31542 20392
rect 31573 20383 31631 20389
rect 31573 20349 31585 20383
rect 31619 20349 31631 20383
rect 31573 20343 31631 20349
rect 26510 20312 26516 20324
rect 26252 20284 26516 20312
rect 23992 20272 23998 20284
rect 26510 20272 26516 20284
rect 26568 20312 26574 20324
rect 27522 20312 27528 20324
rect 26568 20284 27528 20312
rect 26568 20272 26574 20284
rect 27522 20272 27528 20284
rect 27580 20312 27586 20324
rect 31588 20312 31616 20343
rect 32214 20340 32220 20392
rect 32272 20380 32278 20392
rect 32309 20383 32367 20389
rect 32309 20380 32321 20383
rect 32272 20352 32321 20380
rect 32272 20340 32278 20352
rect 32309 20349 32321 20352
rect 32355 20349 32367 20383
rect 32309 20343 32367 20349
rect 32861 20383 32919 20389
rect 32861 20349 32873 20383
rect 32907 20380 32919 20383
rect 33428 20380 33456 20408
rect 32907 20352 33456 20380
rect 35529 20383 35587 20389
rect 32907 20349 32919 20352
rect 32861 20343 32919 20349
rect 35529 20349 35541 20383
rect 35575 20380 35587 20383
rect 35986 20380 35992 20392
rect 35575 20352 35992 20380
rect 35575 20349 35587 20352
rect 35529 20343 35587 20349
rect 32876 20312 32904 20343
rect 35986 20340 35992 20352
rect 36044 20340 36050 20392
rect 38746 20380 38752 20392
rect 38707 20352 38752 20380
rect 38746 20340 38752 20352
rect 38804 20340 38810 20392
rect 40310 20380 40316 20392
rect 40271 20352 40316 20380
rect 40310 20340 40316 20352
rect 40368 20340 40374 20392
rect 44358 20380 44364 20392
rect 44319 20352 44364 20380
rect 44358 20340 44364 20352
rect 44416 20340 44422 20392
rect 44836 20321 44864 20420
rect 45554 20408 45560 20420
rect 45612 20448 45618 20460
rect 45833 20451 45891 20457
rect 45833 20448 45845 20451
rect 45612 20420 45845 20448
rect 45612 20408 45618 20420
rect 45833 20417 45845 20420
rect 45879 20417 45891 20451
rect 45833 20411 45891 20417
rect 46017 20451 46075 20457
rect 46017 20417 46029 20451
rect 46063 20448 46075 20451
rect 46569 20451 46627 20457
rect 46569 20448 46581 20451
rect 46063 20420 46581 20448
rect 46063 20417 46075 20420
rect 46017 20411 46075 20417
rect 46569 20417 46581 20420
rect 46615 20417 46627 20451
rect 46569 20411 46627 20417
rect 48130 20408 48136 20460
rect 48188 20448 48194 20460
rect 48225 20451 48283 20457
rect 48225 20448 48237 20451
rect 48188 20420 48237 20448
rect 48188 20408 48194 20420
rect 48225 20417 48237 20420
rect 48271 20417 48283 20451
rect 48225 20411 48283 20417
rect 48774 20408 48780 20460
rect 48832 20448 48838 20460
rect 49252 20457 49280 20488
rect 49329 20519 49387 20525
rect 49329 20485 49341 20519
rect 49375 20516 49387 20519
rect 49786 20516 49792 20528
rect 49375 20488 49792 20516
rect 49375 20485 49387 20488
rect 49329 20479 49387 20485
rect 49786 20476 49792 20488
rect 49844 20476 49850 20528
rect 50341 20519 50399 20525
rect 50341 20485 50353 20519
rect 50387 20516 50399 20519
rect 50890 20516 50896 20528
rect 50387 20488 50896 20516
rect 50387 20485 50399 20488
rect 50341 20479 50399 20485
rect 50890 20476 50896 20488
rect 50948 20476 50954 20528
rect 51046 20516 51080 20528
rect 51000 20488 51080 20516
rect 48869 20451 48927 20457
rect 48869 20448 48881 20451
rect 48832 20420 48881 20448
rect 48832 20408 48838 20420
rect 48869 20417 48881 20420
rect 48915 20417 48927 20451
rect 48869 20411 48927 20417
rect 48961 20451 49019 20457
rect 48961 20417 48973 20451
rect 49007 20417 49019 20451
rect 48961 20411 49019 20417
rect 49237 20451 49295 20457
rect 49237 20417 49249 20451
rect 49283 20417 49295 20451
rect 50062 20448 50068 20460
rect 50023 20420 50068 20448
rect 49237 20411 49295 20417
rect 45649 20383 45707 20389
rect 45649 20349 45661 20383
rect 45695 20380 45707 20383
rect 45738 20380 45744 20392
rect 45695 20352 45744 20380
rect 45695 20349 45707 20352
rect 45649 20343 45707 20349
rect 45738 20340 45744 20352
rect 45796 20340 45802 20392
rect 48041 20383 48099 20389
rect 48041 20349 48053 20383
rect 48087 20380 48099 20383
rect 48976 20380 49004 20411
rect 50062 20408 50068 20420
rect 50120 20408 50126 20460
rect 50154 20408 50160 20460
rect 50212 20448 50218 20460
rect 51000 20457 51028 20488
rect 51074 20476 51080 20488
rect 51132 20516 51138 20528
rect 51534 20516 51540 20528
rect 51132 20488 51540 20516
rect 51132 20476 51138 20488
rect 51534 20476 51540 20488
rect 51592 20476 51598 20528
rect 51629 20519 51687 20525
rect 51629 20485 51641 20519
rect 51675 20516 51687 20519
rect 54588 20516 54616 20556
rect 55214 20544 55220 20556
rect 55272 20544 55278 20596
rect 56045 20587 56103 20593
rect 56045 20553 56057 20587
rect 56091 20584 56103 20587
rect 57514 20584 57520 20596
rect 56091 20556 57520 20584
rect 56091 20553 56103 20556
rect 56045 20547 56103 20553
rect 57514 20544 57520 20556
rect 57572 20584 57578 20596
rect 58161 20587 58219 20593
rect 58161 20584 58173 20587
rect 57572 20556 58173 20584
rect 57572 20544 57578 20556
rect 58161 20553 58173 20556
rect 58207 20553 58219 20587
rect 58161 20547 58219 20553
rect 54754 20516 54760 20528
rect 51675 20488 54616 20516
rect 54715 20488 54760 20516
rect 51675 20485 51687 20488
rect 51629 20479 51687 20485
rect 54754 20476 54760 20488
rect 54812 20476 54818 20528
rect 56689 20519 56747 20525
rect 56689 20485 56701 20519
rect 56735 20516 56747 20519
rect 56962 20516 56968 20528
rect 56735 20488 56968 20516
rect 56735 20485 56747 20488
rect 56689 20479 56747 20485
rect 56962 20476 56968 20488
rect 57020 20476 57026 20528
rect 57698 20476 57704 20528
rect 57756 20516 57762 20528
rect 58345 20519 58403 20525
rect 58345 20516 58357 20519
rect 57756 20488 58357 20516
rect 57756 20476 57762 20488
rect 58345 20485 58357 20488
rect 58391 20485 58403 20519
rect 58345 20479 58403 20485
rect 50985 20451 51043 20457
rect 50212 20420 50257 20448
rect 50212 20408 50218 20420
rect 50985 20417 50997 20451
rect 51031 20417 51043 20451
rect 51166 20448 51172 20460
rect 51127 20420 51172 20448
rect 50985 20411 51043 20417
rect 51166 20408 51172 20420
rect 51224 20408 51230 20460
rect 51445 20451 51503 20457
rect 51445 20417 51457 20451
rect 51491 20417 51503 20451
rect 51445 20411 51503 20417
rect 48087 20352 49004 20380
rect 50341 20383 50399 20389
rect 48087 20349 48099 20352
rect 48041 20343 48099 20349
rect 48884 20324 48912 20352
rect 50341 20349 50353 20383
rect 50387 20349 50399 20383
rect 50341 20343 50399 20349
rect 27580 20284 32904 20312
rect 44821 20315 44879 20321
rect 27580 20272 27586 20284
rect 44821 20281 44833 20315
rect 44867 20281 44879 20315
rect 44821 20275 44879 20281
rect 48866 20272 48872 20324
rect 48924 20272 48930 20324
rect 50356 20312 50384 20343
rect 50890 20340 50896 20392
rect 50948 20380 50954 20392
rect 51460 20380 51488 20411
rect 52546 20408 52552 20460
rect 52604 20448 52610 20460
rect 52917 20451 52975 20457
rect 52917 20448 52929 20451
rect 52604 20420 52929 20448
rect 52604 20408 52610 20420
rect 52917 20417 52929 20420
rect 52963 20417 52975 20451
rect 54018 20448 54024 20460
rect 52917 20411 52975 20417
rect 53024 20420 54024 20448
rect 50948 20352 51488 20380
rect 50948 20340 50954 20352
rect 52730 20340 52736 20392
rect 52788 20380 52794 20392
rect 53024 20380 53052 20420
rect 54018 20408 54024 20420
rect 54076 20448 54082 20460
rect 54113 20451 54171 20457
rect 54113 20448 54125 20451
rect 54076 20420 54125 20448
rect 54076 20408 54082 20420
rect 54113 20417 54125 20420
rect 54159 20417 54171 20451
rect 54113 20411 54171 20417
rect 54202 20408 54208 20460
rect 54260 20448 54266 20460
rect 54297 20451 54355 20457
rect 54297 20448 54309 20451
rect 54260 20420 54309 20448
rect 54260 20408 54266 20420
rect 54297 20417 54309 20420
rect 54343 20417 54355 20451
rect 54297 20411 54355 20417
rect 54389 20451 54447 20457
rect 54389 20417 54401 20451
rect 54435 20417 54447 20451
rect 54389 20411 54447 20417
rect 53190 20380 53196 20392
rect 52788 20352 53052 20380
rect 53151 20352 53196 20380
rect 52788 20340 52794 20352
rect 53190 20340 53196 20352
rect 53248 20340 53254 20392
rect 54404 20380 54432 20411
rect 54478 20408 54484 20460
rect 54536 20457 54542 20460
rect 54536 20451 54556 20457
rect 54544 20417 54556 20451
rect 54536 20411 54556 20417
rect 54536 20408 54542 20411
rect 55398 20408 55404 20460
rect 55456 20448 55462 20460
rect 55585 20451 55643 20457
rect 55585 20448 55597 20451
rect 55456 20420 55597 20448
rect 55456 20408 55462 20420
rect 55585 20417 55597 20420
rect 55631 20417 55643 20451
rect 56594 20448 56600 20460
rect 56555 20420 56600 20448
rect 55585 20411 55643 20417
rect 56594 20408 56600 20420
rect 56652 20408 56658 20460
rect 56781 20451 56839 20457
rect 56781 20417 56793 20451
rect 56827 20417 56839 20451
rect 56980 20448 57008 20476
rect 58069 20451 58127 20457
rect 58069 20448 58081 20451
rect 56980 20420 58081 20448
rect 56781 20411 56839 20417
rect 58069 20417 58081 20420
rect 58115 20417 58127 20451
rect 58069 20411 58127 20417
rect 54404 20352 54524 20380
rect 53208 20312 53236 20340
rect 54496 20324 54524 20352
rect 56502 20340 56508 20392
rect 56560 20380 56566 20392
rect 56796 20380 56824 20411
rect 56560 20352 56824 20380
rect 56560 20340 56566 20352
rect 50356 20284 53236 20312
rect 54478 20272 54484 20324
rect 54536 20272 54542 20324
rect 58342 20312 58348 20324
rect 58303 20284 58348 20312
rect 58342 20272 58348 20284
rect 58400 20272 58406 20324
rect 36078 20244 36084 20256
rect 36039 20216 36084 20244
rect 36078 20204 36084 20216
rect 36136 20204 36142 20256
rect 36722 20204 36728 20256
rect 36780 20244 36786 20256
rect 36817 20247 36875 20253
rect 36817 20244 36829 20247
rect 36780 20216 36829 20244
rect 36780 20204 36786 20216
rect 36817 20213 36829 20216
rect 36863 20213 36875 20247
rect 36817 20207 36875 20213
rect 41414 20204 41420 20256
rect 41472 20244 41478 20256
rect 41693 20247 41751 20253
rect 41693 20244 41705 20247
rect 41472 20216 41705 20244
rect 41472 20204 41478 20216
rect 41693 20213 41705 20216
rect 41739 20213 41751 20247
rect 42794 20244 42800 20256
rect 42755 20216 42800 20244
rect 41693 20207 41751 20213
rect 42794 20204 42800 20216
rect 42852 20204 42858 20256
rect 49142 20244 49148 20256
rect 49103 20216 49148 20244
rect 49142 20204 49148 20216
rect 49200 20204 49206 20256
rect 51810 20204 51816 20256
rect 51868 20244 51874 20256
rect 52089 20247 52147 20253
rect 52089 20244 52101 20247
rect 51868 20216 52101 20244
rect 51868 20204 51874 20216
rect 52089 20213 52101 20216
rect 52135 20213 52147 20247
rect 53006 20244 53012 20256
rect 52967 20216 53012 20244
rect 52089 20207 52147 20213
rect 53006 20204 53012 20216
rect 53064 20204 53070 20256
rect 54294 20204 54300 20256
rect 54352 20244 54358 20256
rect 54754 20244 54760 20256
rect 54352 20216 54760 20244
rect 54352 20204 54358 20216
rect 54754 20204 54760 20216
rect 54812 20204 54818 20256
rect 55674 20244 55680 20256
rect 55635 20216 55680 20244
rect 55674 20204 55680 20216
rect 55732 20204 55738 20256
rect 56686 20204 56692 20256
rect 56744 20244 56750 20256
rect 57241 20247 57299 20253
rect 57241 20244 57253 20247
rect 56744 20216 57253 20244
rect 56744 20204 56750 20216
rect 57241 20213 57253 20216
rect 57287 20213 57299 20247
rect 57241 20207 57299 20213
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 23477 20043 23535 20049
rect 23477 20009 23489 20043
rect 23523 20040 23535 20043
rect 23566 20040 23572 20052
rect 23523 20012 23572 20040
rect 23523 20009 23535 20012
rect 23477 20003 23535 20009
rect 23566 20000 23572 20012
rect 23624 20000 23630 20052
rect 23934 20040 23940 20052
rect 23895 20012 23940 20040
rect 23934 20000 23940 20012
rect 23992 20000 23998 20052
rect 27062 20040 27068 20052
rect 27023 20012 27068 20040
rect 27062 20000 27068 20012
rect 27120 20000 27126 20052
rect 28258 20000 28264 20052
rect 28316 20040 28322 20052
rect 29730 20040 29736 20052
rect 28316 20012 28994 20040
rect 29691 20012 29736 20040
rect 28316 20000 28322 20012
rect 26510 19972 26516 19984
rect 26471 19944 26516 19972
rect 26510 19932 26516 19944
rect 26568 19932 26574 19984
rect 27982 19932 27988 19984
rect 28040 19972 28046 19984
rect 28626 19972 28632 19984
rect 28040 19944 28632 19972
rect 28040 19932 28046 19944
rect 24486 19864 24492 19916
rect 24544 19904 24550 19916
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 24544 19876 24593 19904
rect 24544 19864 24550 19876
rect 24581 19873 24593 19876
rect 24627 19873 24639 19907
rect 25498 19904 25504 19916
rect 25459 19876 25504 19904
rect 24581 19867 24639 19873
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 28258 19904 28264 19916
rect 26160 19876 26924 19904
rect 28219 19876 28264 19904
rect 23753 19839 23811 19845
rect 23753 19805 23765 19839
rect 23799 19805 23811 19839
rect 24026 19836 24032 19848
rect 23987 19808 24032 19836
rect 23753 19799 23811 19805
rect 23768 19768 23796 19799
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 25314 19836 25320 19848
rect 25275 19808 25320 19836
rect 25314 19796 25320 19808
rect 25372 19836 25378 19848
rect 26160 19836 26188 19876
rect 25372 19808 26188 19836
rect 25372 19796 25378 19808
rect 26234 19796 26240 19848
rect 26292 19836 26298 19848
rect 26418 19836 26424 19848
rect 26292 19808 26424 19836
rect 26292 19796 26298 19808
rect 26418 19796 26424 19808
rect 26476 19836 26482 19848
rect 26789 19839 26847 19845
rect 26789 19836 26801 19839
rect 26476 19808 26801 19836
rect 26476 19796 26482 19808
rect 26789 19805 26801 19808
rect 26835 19805 26847 19839
rect 26896 19836 26924 19876
rect 28258 19864 28264 19876
rect 28316 19864 28322 19916
rect 28460 19913 28488 19944
rect 28626 19932 28632 19944
rect 28684 19932 28690 19984
rect 28445 19907 28503 19913
rect 28445 19873 28457 19907
rect 28491 19873 28503 19907
rect 28966 19904 28994 20012
rect 29730 20000 29736 20012
rect 29788 20000 29794 20052
rect 31573 20043 31631 20049
rect 31573 20009 31585 20043
rect 31619 20040 31631 20043
rect 31662 20040 31668 20052
rect 31619 20012 31668 20040
rect 31619 20009 31631 20012
rect 31573 20003 31631 20009
rect 31662 20000 31668 20012
rect 31720 20000 31726 20052
rect 33502 20040 33508 20052
rect 33463 20012 33508 20040
rect 33502 20000 33508 20012
rect 33560 20000 33566 20052
rect 35253 20043 35311 20049
rect 35253 20009 35265 20043
rect 35299 20040 35311 20043
rect 35434 20040 35440 20052
rect 35299 20012 35440 20040
rect 35299 20009 35311 20012
rect 35253 20003 35311 20009
rect 35434 20000 35440 20012
rect 35492 20000 35498 20052
rect 38105 20043 38163 20049
rect 38105 20009 38117 20043
rect 38151 20040 38163 20043
rect 38838 20040 38844 20052
rect 38151 20012 38844 20040
rect 38151 20009 38163 20012
rect 38105 20003 38163 20009
rect 38838 20000 38844 20012
rect 38896 20000 38902 20052
rect 39022 20000 39028 20052
rect 39080 20040 39086 20052
rect 39209 20043 39267 20049
rect 39209 20040 39221 20043
rect 39080 20012 39221 20040
rect 39080 20000 39086 20012
rect 39209 20009 39221 20012
rect 39255 20009 39267 20043
rect 39209 20003 39267 20009
rect 40405 20043 40463 20049
rect 40405 20009 40417 20043
rect 40451 20040 40463 20043
rect 40586 20040 40592 20052
rect 40451 20012 40592 20040
rect 40451 20009 40463 20012
rect 40405 20003 40463 20009
rect 40586 20000 40592 20012
rect 40644 20000 40650 20052
rect 44358 20040 44364 20052
rect 44319 20012 44364 20040
rect 44358 20000 44364 20012
rect 44416 20000 44422 20052
rect 46937 20043 46995 20049
rect 46937 20009 46949 20043
rect 46983 20040 46995 20043
rect 47118 20040 47124 20052
rect 46983 20012 47124 20040
rect 46983 20009 46995 20012
rect 46937 20003 46995 20009
rect 47118 20000 47124 20012
rect 47176 20000 47182 20052
rect 47394 20040 47400 20052
rect 47355 20012 47400 20040
rect 47394 20000 47400 20012
rect 47452 20000 47458 20052
rect 49142 20040 49148 20052
rect 49103 20012 49148 20040
rect 49142 20000 49148 20012
rect 49200 20000 49206 20052
rect 51166 20000 51172 20052
rect 51224 20040 51230 20052
rect 51629 20043 51687 20049
rect 51629 20040 51641 20043
rect 51224 20012 51641 20040
rect 51224 20000 51230 20012
rect 51629 20009 51641 20012
rect 51675 20009 51687 20043
rect 51629 20003 51687 20009
rect 54202 20000 54208 20052
rect 54260 20040 54266 20052
rect 54481 20043 54539 20049
rect 54481 20040 54493 20043
rect 54260 20012 54493 20040
rect 54260 20000 54266 20012
rect 54481 20009 54493 20012
rect 54527 20009 54539 20043
rect 54481 20003 54539 20009
rect 55769 20043 55827 20049
rect 55769 20009 55781 20043
rect 55815 20040 55827 20043
rect 56318 20040 56324 20052
rect 55815 20012 56324 20040
rect 55815 20009 55827 20012
rect 55769 20003 55827 20009
rect 56318 20000 56324 20012
rect 56376 20000 56382 20052
rect 57698 20000 57704 20052
rect 57756 20040 57762 20052
rect 57793 20043 57851 20049
rect 57793 20040 57805 20043
rect 57756 20012 57805 20040
rect 57756 20000 57762 20012
rect 57793 20009 57805 20012
rect 57839 20009 57851 20043
rect 57793 20003 57851 20009
rect 37185 19975 37243 19981
rect 37185 19941 37197 19975
rect 37231 19972 37243 19975
rect 38746 19972 38752 19984
rect 37231 19944 38752 19972
rect 37231 19941 37243 19944
rect 37185 19935 37243 19941
rect 38746 19932 38752 19944
rect 38804 19932 38810 19984
rect 46290 19932 46296 19984
rect 46348 19972 46354 19984
rect 46569 19975 46627 19981
rect 46569 19972 46581 19975
rect 46348 19944 46581 19972
rect 46348 19932 46354 19944
rect 46569 19941 46581 19944
rect 46615 19972 46627 19975
rect 47673 19975 47731 19981
rect 47673 19972 47685 19975
rect 46615 19944 47685 19972
rect 46615 19941 46627 19944
rect 46569 19935 46627 19941
rect 47673 19941 47685 19944
rect 47719 19941 47731 19975
rect 47673 19935 47731 19941
rect 47762 19932 47768 19984
rect 47820 19972 47826 19984
rect 48590 19972 48596 19984
rect 47820 19944 48596 19972
rect 47820 19932 47826 19944
rect 48590 19932 48596 19944
rect 48648 19932 48654 19984
rect 50893 19975 50951 19981
rect 50893 19941 50905 19975
rect 50939 19972 50951 19975
rect 54018 19972 54024 19984
rect 50939 19944 54024 19972
rect 50939 19941 50951 19944
rect 50893 19935 50951 19941
rect 54018 19932 54024 19944
rect 54076 19932 54082 19984
rect 29270 19904 29276 19916
rect 28966 19876 29276 19904
rect 28445 19867 28503 19873
rect 29270 19864 29276 19876
rect 29328 19864 29334 19916
rect 33410 19904 33416 19916
rect 33323 19876 33416 19904
rect 28350 19836 28356 19848
rect 26896 19808 28356 19836
rect 26789 19799 26847 19805
rect 28350 19796 28356 19808
rect 28408 19796 28414 19848
rect 28530 19839 28588 19845
rect 28530 19805 28542 19839
rect 28576 19805 28588 19839
rect 29914 19836 29920 19848
rect 29875 19808 29920 19836
rect 28530 19799 28588 19805
rect 25038 19768 25044 19780
rect 23768 19740 25044 19768
rect 25038 19728 25044 19740
rect 25096 19728 25102 19780
rect 26602 19728 26608 19780
rect 26660 19768 26666 19780
rect 26881 19771 26939 19777
rect 26881 19768 26893 19771
rect 26660 19740 26893 19768
rect 26660 19728 26666 19740
rect 26881 19737 26893 19740
rect 26927 19737 26939 19771
rect 26881 19731 26939 19737
rect 28552 19712 28580 19799
rect 29914 19796 29920 19808
rect 29972 19796 29978 19848
rect 30009 19839 30067 19845
rect 30009 19805 30021 19839
rect 30055 19805 30067 19839
rect 30009 19799 30067 19805
rect 31481 19839 31539 19845
rect 31481 19805 31493 19839
rect 31527 19836 31539 19839
rect 31570 19836 31576 19848
rect 31527 19808 31576 19836
rect 31527 19805 31539 19808
rect 31481 19799 31539 19805
rect 29546 19728 29552 19780
rect 29604 19768 29610 19780
rect 30024 19768 30052 19799
rect 31570 19796 31576 19808
rect 31628 19796 31634 19848
rect 31665 19839 31723 19845
rect 31665 19805 31677 19839
rect 31711 19836 31723 19839
rect 32214 19836 32220 19848
rect 31711 19808 32220 19836
rect 31711 19805 31723 19808
rect 31665 19799 31723 19805
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 33336 19845 33364 19876
rect 33410 19864 33416 19876
rect 33468 19904 33474 19916
rect 36538 19904 36544 19916
rect 33468 19876 35940 19904
rect 36499 19876 36544 19904
rect 33468 19864 33474 19876
rect 33321 19839 33379 19845
rect 33321 19805 33333 19839
rect 33367 19805 33379 19839
rect 33321 19799 33379 19805
rect 34606 19796 34612 19848
rect 34664 19836 34670 19848
rect 35621 19839 35679 19845
rect 35621 19836 35633 19839
rect 34664 19808 35633 19836
rect 34664 19796 34670 19808
rect 35621 19805 35633 19808
rect 35667 19836 35679 19839
rect 35802 19836 35808 19848
rect 35667 19808 35808 19836
rect 35667 19805 35679 19808
rect 35621 19799 35679 19805
rect 35802 19796 35808 19808
rect 35860 19796 35866 19848
rect 35912 19836 35940 19876
rect 36538 19864 36544 19876
rect 36596 19864 36602 19916
rect 36722 19904 36728 19916
rect 36683 19876 36728 19904
rect 36722 19864 36728 19876
rect 36780 19864 36786 19916
rect 37921 19907 37979 19913
rect 37921 19873 37933 19907
rect 37967 19904 37979 19907
rect 38010 19904 38016 19916
rect 37967 19876 38016 19904
rect 37967 19873 37979 19876
rect 37921 19867 37979 19873
rect 38010 19864 38016 19876
rect 38068 19864 38074 19916
rect 37458 19836 37464 19848
rect 35912 19808 37464 19836
rect 37458 19796 37464 19808
rect 37516 19796 37522 19848
rect 37826 19836 37832 19848
rect 37787 19808 37832 19836
rect 37826 19796 37832 19808
rect 37884 19796 37890 19848
rect 38764 19845 38792 19932
rect 40034 19904 40040 19916
rect 39995 19876 40040 19904
rect 40034 19864 40040 19876
rect 40092 19864 40098 19916
rect 41414 19864 41420 19916
rect 41472 19904 41478 19916
rect 42794 19904 42800 19916
rect 41472 19876 41517 19904
rect 42755 19876 42800 19904
rect 41472 19864 41478 19876
rect 42794 19864 42800 19876
rect 42852 19864 42858 19916
rect 46014 19864 46020 19916
rect 46072 19904 46078 19916
rect 46477 19907 46535 19913
rect 46477 19904 46489 19907
rect 46072 19876 46489 19904
rect 46072 19864 46078 19876
rect 46477 19873 46489 19876
rect 46523 19873 46535 19907
rect 46477 19867 46535 19873
rect 46768 19876 47900 19904
rect 38749 19839 38807 19845
rect 38749 19805 38761 19839
rect 38795 19805 38807 19839
rect 38749 19799 38807 19805
rect 40221 19839 40279 19845
rect 40221 19805 40233 19839
rect 40267 19836 40279 19839
rect 40310 19836 40316 19848
rect 40267 19808 40316 19836
rect 40267 19805 40279 19808
rect 40221 19799 40279 19805
rect 40310 19796 40316 19808
rect 40368 19796 40374 19848
rect 41506 19796 41512 19848
rect 41564 19796 41570 19848
rect 43070 19836 43076 19848
rect 43031 19808 43076 19836
rect 43070 19796 43076 19808
rect 43128 19796 43134 19848
rect 44269 19839 44327 19845
rect 44269 19805 44281 19839
rect 44315 19805 44327 19839
rect 44269 19799 44327 19805
rect 44453 19839 44511 19845
rect 44453 19805 44465 19839
rect 44499 19836 44511 19839
rect 44542 19836 44548 19848
rect 44499 19808 44548 19836
rect 44499 19805 44511 19808
rect 44453 19799 44511 19805
rect 29604 19740 30052 19768
rect 29604 19728 29610 19740
rect 33226 19728 33232 19780
rect 33284 19768 33290 19780
rect 33413 19771 33471 19777
rect 33413 19768 33425 19771
rect 33284 19740 33425 19768
rect 33284 19728 33290 19740
rect 33413 19737 33425 19740
rect 33459 19737 33471 19771
rect 33413 19731 33471 19737
rect 33597 19771 33655 19777
rect 33597 19737 33609 19771
rect 33643 19768 33655 19771
rect 33778 19768 33784 19780
rect 33643 19740 33784 19768
rect 33643 19737 33655 19740
rect 33597 19731 33655 19737
rect 33778 19728 33784 19740
rect 33836 19728 33842 19780
rect 35437 19771 35495 19777
rect 35437 19737 35449 19771
rect 35483 19768 35495 19771
rect 36078 19768 36084 19780
rect 35483 19740 36084 19768
rect 35483 19737 35495 19740
rect 35437 19731 35495 19737
rect 36078 19728 36084 19740
rect 36136 19728 36142 19780
rect 42242 19768 42248 19780
rect 42203 19740 42248 19768
rect 42242 19728 42248 19740
rect 42300 19728 42306 19780
rect 26326 19660 26332 19712
rect 26384 19700 26390 19712
rect 26697 19703 26755 19709
rect 26697 19700 26709 19703
rect 26384 19672 26709 19700
rect 26384 19660 26390 19672
rect 26697 19669 26709 19672
rect 26743 19669 26755 19703
rect 28074 19700 28080 19712
rect 28035 19672 28080 19700
rect 26697 19663 26755 19669
rect 28074 19660 28080 19672
rect 28132 19660 28138 19712
rect 28534 19660 28540 19712
rect 28592 19700 28598 19712
rect 29089 19703 29147 19709
rect 29089 19700 29101 19703
rect 28592 19672 29101 19700
rect 28592 19660 28598 19672
rect 29089 19669 29101 19672
rect 29135 19669 29147 19703
rect 29089 19663 29147 19669
rect 30926 19660 30932 19712
rect 30984 19700 30990 19712
rect 32674 19700 32680 19712
rect 30984 19672 32680 19700
rect 30984 19660 30990 19672
rect 32674 19660 32680 19672
rect 32732 19660 32738 19712
rect 36814 19700 36820 19712
rect 36775 19672 36820 19700
rect 36814 19660 36820 19672
rect 36872 19660 36878 19712
rect 43714 19660 43720 19712
rect 43772 19700 43778 19712
rect 43809 19703 43867 19709
rect 43809 19700 43821 19703
rect 43772 19672 43821 19700
rect 43772 19660 43778 19672
rect 43809 19669 43821 19672
rect 43855 19700 43867 19703
rect 44284 19700 44312 19799
rect 44542 19796 44548 19808
rect 44600 19796 44606 19848
rect 45554 19836 45560 19848
rect 45515 19808 45560 19836
rect 45554 19796 45560 19808
rect 45612 19796 45618 19848
rect 45738 19836 45744 19848
rect 45699 19808 45744 19836
rect 45738 19796 45744 19808
rect 45796 19796 45802 19848
rect 45646 19728 45652 19780
rect 45704 19768 45710 19780
rect 45925 19771 45983 19777
rect 45925 19768 45937 19771
rect 45704 19740 45937 19768
rect 45704 19728 45710 19740
rect 45925 19737 45937 19740
rect 45971 19737 45983 19771
rect 46492 19768 46520 19867
rect 46768 19845 46796 19876
rect 47872 19845 47900 19876
rect 48958 19864 48964 19916
rect 49016 19904 49022 19916
rect 49145 19907 49203 19913
rect 49145 19904 49157 19907
rect 49016 19876 49157 19904
rect 49016 19864 49022 19876
rect 49145 19873 49157 19876
rect 49191 19873 49203 19907
rect 49145 19867 49203 19873
rect 52273 19907 52331 19913
rect 52273 19873 52285 19907
rect 52319 19904 52331 19907
rect 52822 19904 52828 19916
rect 52319 19876 52828 19904
rect 52319 19873 52331 19876
rect 52273 19867 52331 19873
rect 52822 19864 52828 19876
rect 52880 19864 52886 19916
rect 53285 19907 53343 19913
rect 53285 19873 53297 19907
rect 53331 19873 53343 19907
rect 53285 19867 53343 19873
rect 46753 19839 46811 19845
rect 46753 19805 46765 19839
rect 46799 19805 46811 19839
rect 46753 19799 46811 19805
rect 47581 19839 47639 19845
rect 47581 19805 47593 19839
rect 47627 19805 47639 19839
rect 47581 19799 47639 19805
rect 47857 19839 47915 19845
rect 47857 19805 47869 19839
rect 47903 19836 47915 19839
rect 48222 19836 48228 19848
rect 47903 19808 48228 19836
rect 47903 19805 47915 19808
rect 47857 19799 47915 19805
rect 47486 19768 47492 19780
rect 46492 19740 47492 19768
rect 45925 19731 45983 19737
rect 43855 19672 44312 19700
rect 45940 19700 45968 19731
rect 47486 19728 47492 19740
rect 47544 19768 47550 19780
rect 47596 19768 47624 19799
rect 48222 19796 48228 19808
rect 48280 19836 48286 19848
rect 48866 19836 48872 19848
rect 48280 19808 48872 19836
rect 48280 19796 48286 19808
rect 48866 19796 48872 19808
rect 48924 19796 48930 19848
rect 49053 19839 49111 19845
rect 49053 19805 49065 19839
rect 49099 19805 49111 19839
rect 49053 19799 49111 19805
rect 50433 19839 50491 19845
rect 50433 19805 50445 19839
rect 50479 19836 50491 19839
rect 50890 19836 50896 19848
rect 50479 19808 50896 19836
rect 50479 19805 50491 19808
rect 50433 19799 50491 19805
rect 47544 19740 47624 19768
rect 47544 19728 47550 19740
rect 48590 19728 48596 19780
rect 48648 19768 48654 19780
rect 48777 19771 48835 19777
rect 48777 19768 48789 19771
rect 48648 19740 48789 19768
rect 48648 19728 48654 19740
rect 48777 19737 48789 19740
rect 48823 19737 48835 19771
rect 49068 19768 49096 19799
rect 50890 19796 50896 19808
rect 50948 19796 50954 19848
rect 50985 19839 51043 19845
rect 50985 19805 50997 19839
rect 51031 19805 51043 19839
rect 50985 19799 51043 19805
rect 49142 19768 49148 19780
rect 49068 19740 49148 19768
rect 48777 19731 48835 19737
rect 49142 19728 49148 19740
rect 49200 19728 49206 19780
rect 51000 19768 51028 19799
rect 51074 19796 51080 19848
rect 51132 19836 51138 19848
rect 51994 19836 52000 19848
rect 51132 19808 51177 19836
rect 51955 19808 52000 19836
rect 51132 19796 51138 19808
rect 51994 19796 52000 19808
rect 52052 19796 52058 19848
rect 52730 19796 52736 19848
rect 52788 19836 52794 19848
rect 53009 19839 53067 19845
rect 53009 19836 53021 19839
rect 52788 19808 53021 19836
rect 52788 19796 52794 19808
rect 53009 19805 53021 19808
rect 53055 19805 53067 19839
rect 53009 19799 53067 19805
rect 53098 19796 53104 19848
rect 53156 19836 53162 19848
rect 53193 19839 53251 19845
rect 53193 19836 53205 19839
rect 53156 19808 53205 19836
rect 53156 19796 53162 19808
rect 53193 19805 53205 19808
rect 53239 19805 53251 19839
rect 53193 19799 53251 19805
rect 53300 19780 53328 19867
rect 53558 19864 53564 19916
rect 53616 19904 53622 19916
rect 54389 19907 54447 19913
rect 54389 19904 54401 19907
rect 53616 19876 54401 19904
rect 53616 19864 53622 19876
rect 54389 19873 54401 19876
rect 54435 19904 54447 19907
rect 54754 19904 54760 19916
rect 54435 19876 54760 19904
rect 54435 19873 54447 19876
rect 54389 19867 54447 19873
rect 54754 19864 54760 19876
rect 54812 19864 54818 19916
rect 56594 19904 56600 19916
rect 55508 19876 56600 19904
rect 55508 19848 55536 19876
rect 56594 19864 56600 19876
rect 56652 19864 56658 19916
rect 57422 19904 57428 19916
rect 57383 19876 57428 19904
rect 57422 19864 57428 19876
rect 57480 19864 57486 19916
rect 53377 19839 53435 19845
rect 53377 19805 53389 19839
rect 53423 19805 53435 19839
rect 53377 19799 53435 19805
rect 53469 19839 53527 19845
rect 53469 19805 53481 19839
rect 53515 19836 53527 19839
rect 54110 19836 54116 19848
rect 53515 19808 54116 19836
rect 53515 19805 53527 19808
rect 53469 19799 53527 19805
rect 51000 19740 51074 19768
rect 51046 19712 51074 19740
rect 53282 19728 53288 19780
rect 53340 19728 53346 19780
rect 53392 19712 53420 19799
rect 54110 19796 54116 19808
rect 54168 19796 54174 19848
rect 54205 19839 54263 19845
rect 54205 19805 54217 19839
rect 54251 19836 54263 19839
rect 54294 19836 54300 19848
rect 54251 19808 54300 19836
rect 54251 19805 54263 19808
rect 54205 19799 54263 19805
rect 54294 19796 54300 19808
rect 54352 19796 54358 19848
rect 54478 19836 54484 19848
rect 54439 19808 54484 19836
rect 54478 19796 54484 19808
rect 54536 19796 54542 19848
rect 55490 19836 55496 19848
rect 55451 19808 55496 19836
rect 55490 19796 55496 19808
rect 55548 19796 55554 19848
rect 56413 19839 56471 19845
rect 56413 19836 56425 19839
rect 55692 19808 56425 19836
rect 53653 19771 53711 19777
rect 53653 19737 53665 19771
rect 53699 19768 53711 19771
rect 55398 19768 55404 19780
rect 53699 19740 55404 19768
rect 53699 19737 53711 19740
rect 53653 19731 53711 19737
rect 55398 19728 55404 19740
rect 55456 19768 55462 19780
rect 55692 19768 55720 19808
rect 56413 19805 56425 19808
rect 56459 19805 56471 19839
rect 56413 19799 56471 19805
rect 55456 19740 55720 19768
rect 55769 19771 55827 19777
rect 55456 19728 55462 19740
rect 55769 19737 55781 19771
rect 55815 19768 55827 19771
rect 56229 19771 56287 19777
rect 56229 19768 56241 19771
rect 55815 19740 56241 19768
rect 55815 19737 55827 19740
rect 55769 19731 55827 19737
rect 56229 19737 56241 19740
rect 56275 19737 56287 19771
rect 56428 19768 56456 19799
rect 56502 19796 56508 19848
rect 56560 19836 56566 19848
rect 56689 19839 56747 19845
rect 56689 19836 56701 19839
rect 56560 19808 56701 19836
rect 56560 19796 56566 19808
rect 56689 19805 56701 19808
rect 56735 19805 56747 19839
rect 56689 19799 56747 19805
rect 57517 19839 57575 19845
rect 57517 19805 57529 19839
rect 57563 19805 57575 19839
rect 57517 19799 57575 19805
rect 57532 19768 57560 19799
rect 56428 19740 57560 19768
rect 56229 19731 56287 19737
rect 47854 19700 47860 19712
rect 45940 19672 47860 19700
rect 43855 19669 43867 19672
rect 43809 19663 43867 19669
rect 47854 19660 47860 19672
rect 47912 19660 47918 19712
rect 51046 19672 51080 19712
rect 51074 19660 51080 19672
rect 51132 19660 51138 19712
rect 52086 19700 52092 19712
rect 52047 19672 52092 19700
rect 52086 19660 52092 19672
rect 52144 19660 52150 19712
rect 53374 19660 53380 19712
rect 53432 19660 53438 19712
rect 54018 19660 54024 19712
rect 54076 19700 54082 19712
rect 55490 19700 55496 19712
rect 54076 19672 55496 19700
rect 54076 19660 54082 19672
rect 55490 19660 55496 19672
rect 55548 19660 55554 19712
rect 55585 19703 55643 19709
rect 55585 19669 55597 19703
rect 55631 19700 55643 19703
rect 56410 19700 56416 19712
rect 55631 19672 56416 19700
rect 55631 19669 55643 19672
rect 55585 19663 55643 19669
rect 56410 19660 56416 19672
rect 56468 19660 56474 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 23750 19496 23756 19508
rect 23663 19468 23756 19496
rect 23750 19456 23756 19468
rect 23808 19496 23814 19508
rect 24673 19499 24731 19505
rect 23808 19468 24440 19496
rect 23808 19456 23814 19468
rect 24412 19369 24440 19468
rect 24673 19465 24685 19499
rect 24719 19496 24731 19499
rect 25038 19496 25044 19508
rect 24719 19468 25044 19496
rect 24719 19465 24731 19468
rect 24673 19459 24731 19465
rect 25038 19456 25044 19468
rect 25096 19456 25102 19508
rect 25498 19496 25504 19508
rect 25459 19468 25504 19496
rect 25498 19456 25504 19468
rect 25556 19456 25562 19508
rect 26050 19496 26056 19508
rect 26011 19468 26056 19496
rect 26050 19456 26056 19468
rect 26108 19456 26114 19508
rect 34606 19496 34612 19508
rect 29564 19468 34612 19496
rect 28626 19428 28632 19440
rect 25608 19400 28632 19428
rect 24397 19363 24455 19369
rect 22005 19295 22063 19301
rect 22005 19261 22017 19295
rect 22051 19261 22063 19295
rect 22278 19292 22284 19304
rect 22239 19264 22284 19292
rect 22005 19255 22063 19261
rect 22020 19156 22048 19255
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 23400 19292 23428 19346
rect 24397 19329 24409 19363
rect 24443 19329 24455 19363
rect 24397 19323 24455 19329
rect 24765 19363 24823 19369
rect 24765 19329 24777 19363
rect 24811 19329 24823 19363
rect 25406 19360 25412 19372
rect 25367 19332 25412 19360
rect 24765 19323 24823 19329
rect 23842 19292 23848 19304
rect 23400 19264 23848 19292
rect 23842 19252 23848 19264
rect 23900 19252 23906 19304
rect 24780 19292 24808 19323
rect 25406 19320 25412 19332
rect 25464 19320 25470 19372
rect 25608 19369 25636 19400
rect 28626 19388 28632 19400
rect 28684 19388 28690 19440
rect 29564 19437 29592 19468
rect 34606 19456 34612 19468
rect 34664 19456 34670 19508
rect 34698 19456 34704 19508
rect 34756 19496 34762 19508
rect 34885 19499 34943 19505
rect 34885 19496 34897 19499
rect 34756 19468 34897 19496
rect 34756 19456 34762 19468
rect 34885 19465 34897 19468
rect 34931 19465 34943 19499
rect 36906 19496 36912 19508
rect 36867 19468 36912 19496
rect 34885 19459 34943 19465
rect 36906 19456 36912 19468
rect 36964 19456 36970 19508
rect 37921 19499 37979 19505
rect 37921 19465 37933 19499
rect 37967 19496 37979 19499
rect 39114 19496 39120 19508
rect 37967 19468 39120 19496
rect 37967 19465 37979 19468
rect 37921 19459 37979 19465
rect 39114 19456 39120 19468
rect 39172 19456 39178 19508
rect 41230 19496 41236 19508
rect 41191 19468 41236 19496
rect 41230 19456 41236 19468
rect 41288 19456 41294 19508
rect 41874 19496 41880 19508
rect 41835 19468 41880 19496
rect 41874 19456 41880 19468
rect 41932 19456 41938 19508
rect 42797 19499 42855 19505
rect 42797 19465 42809 19499
rect 42843 19496 42855 19499
rect 43070 19496 43076 19508
rect 42843 19468 43076 19496
rect 42843 19465 42855 19468
rect 42797 19459 42855 19465
rect 43070 19456 43076 19468
rect 43128 19456 43134 19508
rect 43714 19496 43720 19508
rect 43675 19468 43720 19496
rect 43714 19456 43720 19468
rect 43772 19456 43778 19508
rect 48133 19499 48191 19505
rect 48133 19465 48145 19499
rect 48179 19496 48191 19499
rect 48222 19496 48228 19508
rect 48179 19468 48228 19496
rect 48179 19465 48191 19468
rect 48133 19459 48191 19465
rect 48222 19456 48228 19468
rect 48280 19456 48286 19508
rect 48590 19456 48596 19508
rect 48648 19496 48654 19508
rect 48648 19468 49096 19496
rect 48648 19456 48654 19468
rect 28813 19431 28871 19437
rect 28813 19397 28825 19431
rect 28859 19428 28871 19431
rect 29549 19431 29607 19437
rect 28859 19400 29500 19428
rect 28859 19397 28871 19400
rect 28813 19391 28871 19397
rect 25593 19363 25651 19369
rect 25593 19329 25605 19363
rect 25639 19329 25651 19363
rect 25593 19323 25651 19329
rect 26421 19363 26479 19369
rect 26421 19329 26433 19363
rect 26467 19360 26479 19363
rect 28074 19360 28080 19372
rect 26467 19332 26740 19360
rect 28035 19332 28080 19360
rect 26467 19329 26479 19332
rect 26421 19323 26479 19329
rect 26234 19292 26240 19304
rect 24780 19264 25176 19292
rect 26195 19264 26240 19292
rect 25148 19236 25176 19264
rect 26234 19252 26240 19264
rect 26292 19252 26298 19304
rect 26326 19252 26332 19304
rect 26384 19292 26390 19304
rect 26384 19264 26429 19292
rect 26384 19252 26390 19264
rect 26510 19252 26516 19304
rect 26568 19292 26574 19304
rect 26712 19292 26740 19332
rect 28074 19320 28080 19332
rect 28132 19320 28138 19372
rect 28350 19320 28356 19372
rect 28408 19360 28414 19372
rect 28721 19363 28779 19369
rect 28721 19360 28733 19363
rect 28408 19332 28733 19360
rect 28408 19320 28414 19332
rect 28721 19329 28733 19332
rect 28767 19329 28779 19363
rect 28902 19360 28908 19372
rect 28863 19332 28908 19360
rect 28721 19323 28779 19329
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29472 19360 29500 19400
rect 29549 19397 29561 19431
rect 29595 19397 29607 19431
rect 29549 19391 29607 19397
rect 32674 19388 32680 19440
rect 32732 19428 32738 19440
rect 33597 19431 33655 19437
rect 33597 19428 33609 19431
rect 32732 19400 33609 19428
rect 32732 19388 32738 19400
rect 33597 19397 33609 19400
rect 33643 19397 33655 19431
rect 34514 19428 34520 19440
rect 33597 19391 33655 19397
rect 34256 19400 34520 19428
rect 29914 19360 29920 19372
rect 29472 19332 29920 19360
rect 29914 19320 29920 19332
rect 29972 19320 29978 19372
rect 30009 19363 30067 19369
rect 30009 19329 30021 19363
rect 30055 19360 30067 19363
rect 30374 19360 30380 19372
rect 30055 19332 30380 19360
rect 30055 19329 30067 19332
rect 30009 19323 30067 19329
rect 30374 19320 30380 19332
rect 30432 19320 30438 19372
rect 31570 19360 31576 19372
rect 31531 19332 31576 19360
rect 31570 19320 31576 19332
rect 31628 19320 31634 19372
rect 31757 19363 31815 19369
rect 31757 19329 31769 19363
rect 31803 19360 31815 19363
rect 32214 19360 32220 19372
rect 31803 19332 32220 19360
rect 31803 19329 31815 19332
rect 31757 19323 31815 19329
rect 32214 19320 32220 19332
rect 32272 19320 32278 19372
rect 32398 19320 32404 19372
rect 32456 19360 32462 19372
rect 32585 19363 32643 19369
rect 32585 19360 32597 19363
rect 32456 19332 32597 19360
rect 32456 19320 32462 19332
rect 32585 19329 32597 19332
rect 32631 19329 32643 19363
rect 32585 19323 32643 19329
rect 33134 19320 33140 19372
rect 33192 19360 33198 19372
rect 34256 19369 34284 19400
rect 34514 19388 34520 19400
rect 34572 19388 34578 19440
rect 36354 19388 36360 19440
rect 36412 19428 36418 19440
rect 36449 19431 36507 19437
rect 36449 19428 36461 19431
rect 36412 19400 36461 19428
rect 36412 19388 36418 19400
rect 36449 19397 36461 19400
rect 36495 19397 36507 19431
rect 39390 19428 39396 19440
rect 39303 19400 39396 19428
rect 36449 19391 36507 19397
rect 39390 19388 39396 19400
rect 39448 19428 39454 19440
rect 39850 19428 39856 19440
rect 39448 19400 39856 19428
rect 39448 19388 39454 19400
rect 39850 19388 39856 19400
rect 39908 19388 39914 19440
rect 40034 19388 40040 19440
rect 40092 19437 40098 19440
rect 40092 19431 40111 19437
rect 40099 19397 40111 19431
rect 40092 19391 40111 19397
rect 40092 19388 40098 19391
rect 45738 19388 45744 19440
rect 45796 19428 45802 19440
rect 46661 19431 46719 19437
rect 46661 19428 46673 19431
rect 45796 19400 46673 19428
rect 45796 19388 45802 19400
rect 46661 19397 46673 19400
rect 46707 19397 46719 19431
rect 48240 19428 48268 19456
rect 48240 19400 48820 19428
rect 46661 19391 46719 19397
rect 33413 19363 33471 19369
rect 33413 19360 33425 19363
rect 33192 19332 33425 19360
rect 33192 19320 33198 19332
rect 33413 19329 33425 19332
rect 33459 19329 33471 19363
rect 33413 19323 33471 19329
rect 34241 19363 34299 19369
rect 34241 19329 34253 19363
rect 34287 19329 34299 19363
rect 34422 19360 34428 19372
rect 34383 19332 34428 19360
rect 34241 19323 34299 19329
rect 34422 19320 34428 19332
rect 34480 19320 34486 19372
rect 34701 19369 34759 19375
rect 34701 19335 34713 19369
rect 34747 19335 34759 19369
rect 34701 19329 34759 19335
rect 27154 19292 27160 19304
rect 26568 19264 26613 19292
rect 26712 19264 27160 19292
rect 26568 19252 26574 19264
rect 25130 19184 25136 19236
rect 25188 19224 25194 19236
rect 26712 19224 26740 19264
rect 27154 19252 27160 19264
rect 27212 19252 27218 19304
rect 27706 19292 27712 19304
rect 27667 19264 27712 19292
rect 27706 19252 27712 19264
rect 27764 19252 27770 19304
rect 28169 19295 28227 19301
rect 28169 19261 28181 19295
rect 28215 19292 28227 19295
rect 29638 19292 29644 19304
rect 28215 19264 29644 19292
rect 28215 19261 28227 19264
rect 28169 19255 28227 19261
rect 29638 19252 29644 19264
rect 29696 19292 29702 19304
rect 29733 19295 29791 19301
rect 29733 19292 29745 19295
rect 29696 19264 29745 19292
rect 29696 19252 29702 19264
rect 29733 19261 29745 19264
rect 29779 19261 29791 19295
rect 29733 19255 29791 19261
rect 29822 19252 29828 19304
rect 29880 19292 29886 19304
rect 31846 19292 31852 19304
rect 29880 19264 29925 19292
rect 30484 19264 31852 19292
rect 29880 19252 29886 19264
rect 25188 19196 26740 19224
rect 25188 19184 25194 19196
rect 29546 19184 29552 19236
rect 29604 19224 29610 19236
rect 30484 19224 30512 19264
rect 31846 19252 31852 19264
rect 31904 19292 31910 19304
rect 32490 19292 32496 19304
rect 31904 19264 32352 19292
rect 32451 19264 32496 19292
rect 31904 19252 31910 19264
rect 29604 19196 30512 19224
rect 31389 19227 31447 19233
rect 29604 19184 29610 19196
rect 31389 19193 31401 19227
rect 31435 19224 31447 19227
rect 31754 19224 31760 19236
rect 31435 19196 31760 19224
rect 31435 19193 31447 19196
rect 31389 19187 31447 19193
rect 31754 19184 31760 19196
rect 31812 19184 31818 19236
rect 32324 19224 32352 19264
rect 32490 19252 32496 19264
rect 32548 19252 32554 19304
rect 32953 19295 33011 19301
rect 32953 19261 32965 19295
rect 32999 19292 33011 19295
rect 33226 19292 33232 19304
rect 32999 19264 33232 19292
rect 32999 19261 33011 19264
rect 32953 19255 33011 19261
rect 33226 19252 33232 19264
rect 33284 19252 33290 19304
rect 33781 19295 33839 19301
rect 33781 19261 33793 19295
rect 33827 19292 33839 19295
rect 34716 19292 34744 19329
rect 34882 19320 34888 19372
rect 34940 19360 34946 19372
rect 35345 19363 35403 19369
rect 35345 19360 35357 19363
rect 34940 19332 35357 19360
rect 34940 19320 34946 19332
rect 35345 19329 35357 19332
rect 35391 19329 35403 19363
rect 35526 19360 35532 19372
rect 35487 19332 35532 19360
rect 35345 19323 35403 19329
rect 35526 19320 35532 19332
rect 35584 19320 35590 19372
rect 35805 19363 35863 19369
rect 35805 19329 35817 19363
rect 35851 19360 35863 19363
rect 35989 19363 36047 19369
rect 35851 19332 35885 19360
rect 35851 19329 35863 19332
rect 35805 19323 35863 19329
rect 35989 19329 36001 19363
rect 36035 19360 36047 19363
rect 37826 19360 37832 19372
rect 36035 19332 37832 19360
rect 36035 19329 36047 19332
rect 35989 19323 36047 19329
rect 34790 19292 34796 19304
rect 33827 19264 34796 19292
rect 33827 19261 33839 19264
rect 33781 19255 33839 19261
rect 34790 19252 34796 19264
rect 34848 19292 34854 19304
rect 35820 19292 35848 19323
rect 37826 19320 37832 19332
rect 37884 19320 37890 19372
rect 38010 19360 38016 19372
rect 37971 19332 38016 19360
rect 38010 19320 38016 19332
rect 38068 19320 38074 19372
rect 41138 19360 41144 19372
rect 41099 19332 41144 19360
rect 41138 19320 41144 19332
rect 41196 19320 41202 19372
rect 41414 19320 41420 19372
rect 41472 19360 41478 19372
rect 41785 19363 41843 19369
rect 41785 19360 41797 19363
rect 41472 19332 41797 19360
rect 41472 19320 41478 19332
rect 41785 19329 41797 19332
rect 41831 19329 41843 19363
rect 41785 19323 41843 19329
rect 41874 19320 41880 19372
rect 41932 19360 41938 19372
rect 41969 19363 42027 19369
rect 41969 19360 41981 19363
rect 41932 19332 41981 19360
rect 41932 19320 41938 19332
rect 41969 19329 41981 19332
rect 42015 19329 42027 19363
rect 41969 19323 42027 19329
rect 42613 19363 42671 19369
rect 42613 19329 42625 19363
rect 42659 19360 42671 19363
rect 42794 19360 42800 19372
rect 42659 19332 42800 19360
rect 42659 19329 42671 19332
rect 42613 19323 42671 19329
rect 42794 19320 42800 19332
rect 42852 19320 42858 19372
rect 43622 19360 43628 19372
rect 43583 19332 43628 19360
rect 43622 19320 43628 19332
rect 43680 19360 43686 19372
rect 44082 19360 44088 19372
rect 43680 19332 44088 19360
rect 43680 19320 43686 19332
rect 44082 19320 44088 19332
rect 44140 19360 44146 19372
rect 46014 19360 46020 19372
rect 44140 19332 45048 19360
rect 45975 19332 46020 19360
rect 44140 19320 44146 19332
rect 45020 19304 45048 19332
rect 46014 19320 46020 19332
rect 46072 19320 46078 19372
rect 48792 19369 48820 19400
rect 49068 19369 49096 19468
rect 50154 19456 50160 19508
rect 50212 19496 50218 19508
rect 50617 19499 50675 19505
rect 50617 19496 50629 19499
rect 50212 19468 50629 19496
rect 50212 19456 50218 19468
rect 50617 19465 50629 19468
rect 50663 19465 50675 19499
rect 51350 19496 51356 19508
rect 51311 19468 51356 19496
rect 50617 19459 50675 19465
rect 51350 19456 51356 19468
rect 51408 19456 51414 19508
rect 51721 19499 51779 19505
rect 51721 19465 51733 19499
rect 51767 19496 51779 19499
rect 52086 19496 52092 19508
rect 51767 19468 52092 19496
rect 51767 19465 51779 19468
rect 51721 19459 51779 19465
rect 52086 19456 52092 19468
rect 52144 19456 52150 19508
rect 53098 19496 53104 19508
rect 53059 19468 53104 19496
rect 53098 19456 53104 19468
rect 53156 19456 53162 19508
rect 54938 19456 54944 19508
rect 54996 19496 55002 19508
rect 55107 19499 55165 19505
rect 55107 19496 55119 19499
rect 54996 19468 55119 19496
rect 54996 19456 55002 19468
rect 55107 19465 55119 19468
rect 55153 19465 55165 19499
rect 55107 19459 55165 19465
rect 57149 19499 57207 19505
rect 57149 19465 57161 19499
rect 57195 19496 57207 19499
rect 57422 19496 57428 19508
rect 57195 19468 57428 19496
rect 57195 19465 57207 19468
rect 57149 19459 57207 19465
rect 57422 19456 57428 19468
rect 57480 19456 57486 19508
rect 51813 19431 51871 19437
rect 51813 19428 51825 19431
rect 50172 19400 51825 19428
rect 50172 19372 50200 19400
rect 51813 19397 51825 19400
rect 51859 19428 51871 19431
rect 51994 19428 52000 19440
rect 51859 19400 52000 19428
rect 51859 19397 51871 19400
rect 51813 19391 51871 19397
rect 51994 19388 52000 19400
rect 52052 19388 52058 19440
rect 48225 19363 48283 19369
rect 48225 19360 48237 19363
rect 47504 19332 48237 19360
rect 34848 19264 35848 19292
rect 43901 19295 43959 19301
rect 34848 19252 34854 19264
rect 43901 19261 43913 19295
rect 43947 19292 43959 19295
rect 43990 19292 43996 19304
rect 43947 19264 43996 19292
rect 43947 19261 43959 19264
rect 43901 19255 43959 19261
rect 43990 19252 43996 19264
rect 44048 19292 44054 19304
rect 44453 19295 44511 19301
rect 44453 19292 44465 19295
rect 44048 19264 44465 19292
rect 44048 19252 44054 19264
rect 44453 19261 44465 19264
rect 44499 19292 44511 19295
rect 44542 19292 44548 19304
rect 44499 19264 44548 19292
rect 44499 19261 44511 19264
rect 44453 19255 44511 19261
rect 44542 19252 44548 19264
rect 44600 19252 44606 19304
rect 45002 19292 45008 19304
rect 44915 19264 45008 19292
rect 45002 19252 45008 19264
rect 45060 19252 45066 19304
rect 46109 19295 46167 19301
rect 46109 19261 46121 19295
rect 46155 19292 46167 19295
rect 46290 19292 46296 19304
rect 46155 19264 46296 19292
rect 46155 19261 46167 19264
rect 46109 19255 46167 19261
rect 46290 19252 46296 19264
rect 46348 19252 46354 19304
rect 46750 19252 46756 19304
rect 46808 19292 46814 19304
rect 47504 19292 47532 19332
rect 46808 19264 47532 19292
rect 46808 19252 46814 19264
rect 36538 19224 36544 19236
rect 32324 19196 36544 19224
rect 36538 19184 36544 19196
rect 36596 19184 36602 19236
rect 36722 19224 36728 19236
rect 36683 19196 36728 19224
rect 36722 19184 36728 19196
rect 36780 19184 36786 19236
rect 22094 19156 22100 19168
rect 22020 19128 22100 19156
rect 22094 19116 22100 19128
rect 22152 19116 22158 19168
rect 25406 19116 25412 19168
rect 25464 19156 25470 19168
rect 27157 19159 27215 19165
rect 27157 19156 27169 19159
rect 25464 19128 27169 19156
rect 25464 19116 25470 19128
rect 27157 19125 27169 19128
rect 27203 19156 27215 19159
rect 28534 19156 28540 19168
rect 27203 19128 28540 19156
rect 27203 19125 27215 19128
rect 27157 19119 27215 19125
rect 28534 19116 28540 19128
rect 28592 19116 28598 19168
rect 40034 19156 40040 19168
rect 39995 19128 40040 19156
rect 40034 19116 40040 19128
rect 40092 19116 40098 19168
rect 40218 19156 40224 19168
rect 40179 19128 40224 19156
rect 40218 19116 40224 19128
rect 40276 19116 40282 19168
rect 43254 19156 43260 19168
rect 43215 19128 43260 19156
rect 43254 19116 43260 19128
rect 43312 19116 43318 19168
rect 45741 19159 45799 19165
rect 45741 19125 45753 19159
rect 45787 19156 45799 19159
rect 45830 19156 45836 19168
rect 45787 19128 45836 19156
rect 45787 19125 45799 19128
rect 45741 19119 45799 19125
rect 45830 19116 45836 19128
rect 45888 19116 45894 19168
rect 48056 19156 48084 19332
rect 48225 19329 48237 19332
rect 48271 19329 48283 19363
rect 48225 19323 48283 19329
rect 48777 19363 48835 19369
rect 48777 19329 48789 19363
rect 48823 19329 48835 19363
rect 48777 19323 48835 19329
rect 49053 19363 49111 19369
rect 49053 19329 49065 19363
rect 49099 19329 49111 19363
rect 49053 19323 49111 19329
rect 49329 19363 49387 19369
rect 49329 19329 49341 19363
rect 49375 19360 49387 19363
rect 50154 19360 50160 19372
rect 49375 19332 50160 19360
rect 49375 19329 49387 19332
rect 49329 19323 49387 19329
rect 50154 19320 50160 19332
rect 50212 19320 50218 19372
rect 50249 19363 50307 19369
rect 50249 19329 50261 19363
rect 50295 19360 50307 19363
rect 52104 19360 52132 19456
rect 55585 19431 55643 19437
rect 55585 19397 55597 19431
rect 55631 19428 55643 19431
rect 56042 19428 56048 19440
rect 55631 19400 56048 19428
rect 55631 19397 55643 19400
rect 55585 19391 55643 19397
rect 56042 19388 56048 19400
rect 56100 19388 56106 19440
rect 53374 19360 53380 19372
rect 50295 19332 52132 19360
rect 53335 19332 53380 19360
rect 50295 19329 50307 19332
rect 50249 19323 50307 19329
rect 48130 19252 48136 19304
rect 48188 19292 48194 19304
rect 48957 19295 49015 19301
rect 48957 19292 48969 19295
rect 48188 19264 48969 19292
rect 48188 19252 48194 19264
rect 48957 19261 48969 19264
rect 49003 19261 49015 19295
rect 49970 19292 49976 19304
rect 49931 19264 49976 19292
rect 48957 19255 49015 19261
rect 49970 19252 49976 19264
rect 50028 19252 50034 19304
rect 50264 19292 50292 19323
rect 53374 19320 53380 19332
rect 53432 19360 53438 19372
rect 54110 19360 54116 19372
rect 53432 19332 54116 19360
rect 53432 19320 53438 19332
rect 54110 19320 54116 19332
rect 54168 19320 54174 19372
rect 56410 19320 56416 19372
rect 56468 19360 56474 19372
rect 56781 19363 56839 19369
rect 56781 19360 56793 19363
rect 56468 19332 56793 19360
rect 56468 19320 56474 19332
rect 56781 19329 56793 19332
rect 56827 19329 56839 19363
rect 56781 19323 56839 19329
rect 51994 19292 52000 19304
rect 50172 19264 50292 19292
rect 51955 19264 52000 19292
rect 48774 19184 48780 19236
rect 48832 19224 48838 19236
rect 48869 19227 48927 19233
rect 48869 19224 48881 19227
rect 48832 19196 48881 19224
rect 48832 19184 48838 19196
rect 48869 19193 48881 19196
rect 48915 19224 48927 19227
rect 49142 19224 49148 19236
rect 48915 19196 49148 19224
rect 48915 19193 48927 19196
rect 48869 19187 48927 19193
rect 49142 19184 49148 19196
rect 49200 19184 49206 19236
rect 50172 19156 50200 19264
rect 51994 19252 52000 19264
rect 52052 19252 52058 19304
rect 53101 19295 53159 19301
rect 53101 19261 53113 19295
rect 53147 19292 53159 19295
rect 53558 19292 53564 19304
rect 53147 19264 53564 19292
rect 53147 19261 53159 19264
rect 53101 19255 53159 19261
rect 53558 19252 53564 19264
rect 53616 19252 53622 19304
rect 55490 19292 55496 19304
rect 55451 19264 55496 19292
rect 55490 19252 55496 19264
rect 55548 19252 55554 19304
rect 55677 19295 55735 19301
rect 55677 19261 55689 19295
rect 55723 19292 55735 19295
rect 55950 19292 55956 19304
rect 55723 19264 55956 19292
rect 55723 19261 55735 19264
rect 55677 19255 55735 19261
rect 55950 19252 55956 19264
rect 56008 19252 56014 19304
rect 56594 19252 56600 19304
rect 56652 19292 56658 19304
rect 56689 19295 56747 19301
rect 56689 19292 56701 19295
rect 56652 19264 56701 19292
rect 56652 19252 56658 19264
rect 56689 19261 56701 19264
rect 56735 19261 56747 19295
rect 56689 19255 56747 19261
rect 50706 19156 50712 19168
rect 48056 19128 50712 19156
rect 50706 19116 50712 19128
rect 50764 19116 50770 19168
rect 53282 19156 53288 19168
rect 53243 19128 53288 19156
rect 53282 19116 53288 19128
rect 53340 19116 53346 19168
rect 53650 19116 53656 19168
rect 53708 19156 53714 19168
rect 53837 19159 53895 19165
rect 53837 19156 53849 19159
rect 53708 19128 53849 19156
rect 53708 19116 53714 19128
rect 53837 19125 53849 19128
rect 53883 19156 53895 19159
rect 54389 19159 54447 19165
rect 54389 19156 54401 19159
rect 53883 19128 54401 19156
rect 53883 19125 53895 19128
rect 53837 19119 53895 19125
rect 54389 19125 54401 19128
rect 54435 19125 54447 19159
rect 54389 19119 54447 19125
rect 58161 19159 58219 19165
rect 58161 19125 58173 19159
rect 58207 19156 58219 19159
rect 58342 19156 58348 19168
rect 58207 19128 58348 19156
rect 58207 19125 58219 19128
rect 58161 19119 58219 19125
rect 58342 19116 58348 19128
rect 58400 19116 58406 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 22097 18955 22155 18961
rect 22097 18921 22109 18955
rect 22143 18952 22155 18955
rect 22278 18952 22284 18964
rect 22143 18924 22284 18952
rect 22143 18921 22155 18924
rect 22097 18915 22155 18921
rect 22278 18912 22284 18924
rect 22336 18912 22342 18964
rect 23845 18955 23903 18961
rect 23845 18921 23857 18955
rect 23891 18952 23903 18955
rect 27522 18952 27528 18964
rect 23891 18924 27528 18952
rect 23891 18921 23903 18924
rect 23845 18915 23903 18921
rect 23860 18816 23888 18915
rect 27522 18912 27528 18924
rect 27580 18912 27586 18964
rect 29089 18955 29147 18961
rect 29089 18921 29101 18955
rect 29135 18952 29147 18955
rect 29822 18952 29828 18964
rect 29135 18924 29828 18952
rect 29135 18921 29147 18924
rect 29089 18915 29147 18921
rect 29822 18912 29828 18924
rect 29880 18912 29886 18964
rect 30558 18912 30564 18964
rect 30616 18952 30622 18964
rect 30745 18955 30803 18961
rect 30745 18952 30757 18955
rect 30616 18924 30757 18952
rect 30616 18912 30622 18924
rect 30745 18921 30757 18924
rect 30791 18921 30803 18955
rect 31570 18952 31576 18964
rect 31531 18924 31576 18952
rect 30745 18915 30803 18921
rect 31570 18912 31576 18924
rect 31628 18912 31634 18964
rect 32490 18952 32496 18964
rect 32451 18924 32496 18952
rect 32490 18912 32496 18924
rect 32548 18912 32554 18964
rect 34790 18912 34796 18964
rect 34848 18952 34854 18964
rect 34885 18955 34943 18961
rect 34885 18952 34897 18955
rect 34848 18924 34897 18952
rect 34848 18912 34854 18924
rect 34885 18921 34897 18924
rect 34931 18921 34943 18955
rect 34885 18915 34943 18921
rect 35161 18955 35219 18961
rect 35161 18921 35173 18955
rect 35207 18952 35219 18955
rect 35618 18952 35624 18964
rect 35207 18924 35624 18952
rect 35207 18921 35219 18924
rect 35161 18915 35219 18921
rect 35618 18912 35624 18924
rect 35676 18912 35682 18964
rect 37550 18912 37556 18964
rect 37608 18952 37614 18964
rect 38197 18955 38255 18961
rect 38197 18952 38209 18955
rect 37608 18924 38209 18952
rect 37608 18912 37614 18924
rect 38197 18921 38209 18924
rect 38243 18921 38255 18955
rect 38197 18915 38255 18921
rect 39209 18955 39267 18961
rect 39209 18921 39221 18955
rect 39255 18952 39267 18955
rect 40034 18952 40040 18964
rect 39255 18924 40040 18952
rect 39255 18921 39267 18924
rect 39209 18915 39267 18921
rect 40034 18912 40040 18924
rect 40092 18912 40098 18964
rect 40310 18912 40316 18964
rect 40368 18952 40374 18964
rect 40773 18955 40831 18961
rect 40773 18952 40785 18955
rect 40368 18924 40785 18952
rect 40368 18912 40374 18924
rect 40773 18921 40785 18924
rect 40819 18921 40831 18955
rect 42794 18952 42800 18964
rect 42755 18924 42800 18952
rect 40773 18915 40831 18921
rect 42794 18912 42800 18924
rect 42852 18912 42858 18964
rect 46014 18912 46020 18964
rect 46072 18952 46078 18964
rect 46477 18955 46535 18961
rect 46477 18952 46489 18955
rect 46072 18924 46489 18952
rect 46072 18912 46078 18924
rect 46477 18921 46489 18924
rect 46523 18921 46535 18955
rect 47486 18952 47492 18964
rect 47447 18924 47492 18952
rect 46477 18915 46535 18921
rect 47486 18912 47492 18924
rect 47544 18912 47550 18964
rect 51074 18912 51080 18964
rect 51132 18952 51138 18964
rect 55490 18952 55496 18964
rect 51132 18924 51177 18952
rect 55451 18924 55496 18952
rect 51132 18912 51138 18924
rect 55490 18912 55496 18924
rect 55548 18912 55554 18964
rect 26605 18887 26663 18893
rect 26605 18853 26617 18887
rect 26651 18884 26663 18887
rect 26694 18884 26700 18896
rect 26651 18856 26700 18884
rect 26651 18853 26663 18856
rect 26605 18847 26663 18853
rect 26694 18844 26700 18856
rect 26752 18844 26758 18896
rect 36924 18856 38976 18884
rect 23124 18788 23888 18816
rect 23124 18757 23152 18788
rect 30006 18776 30012 18828
rect 30064 18816 30070 18828
rect 30285 18819 30343 18825
rect 30285 18816 30297 18819
rect 30064 18788 30297 18816
rect 30064 18776 30070 18788
rect 30285 18785 30297 18788
rect 30331 18785 30343 18819
rect 32769 18819 32827 18825
rect 32769 18816 32781 18819
rect 30285 18779 30343 18785
rect 32140 18788 32781 18816
rect 32140 18760 32168 18788
rect 32769 18785 32781 18788
rect 32815 18785 32827 18819
rect 32769 18779 32827 18785
rect 32861 18819 32919 18825
rect 32861 18785 32873 18819
rect 32907 18816 32919 18819
rect 33226 18816 33232 18828
rect 32907 18788 33232 18816
rect 32907 18785 32919 18788
rect 32861 18779 32919 18785
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18748 21603 18751
rect 22005 18751 22063 18757
rect 22005 18748 22017 18751
rect 21591 18720 22017 18748
rect 21591 18717 21603 18720
rect 21545 18711 21603 18717
rect 22005 18717 22017 18720
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 22189 18751 22247 18757
rect 22189 18717 22201 18751
rect 22235 18717 22247 18751
rect 22189 18711 22247 18717
rect 23109 18751 23167 18757
rect 23109 18717 23121 18751
rect 23155 18717 23167 18751
rect 23109 18711 23167 18717
rect 23293 18751 23351 18757
rect 23293 18717 23305 18751
rect 23339 18748 23351 18751
rect 23750 18748 23756 18760
rect 23339 18720 23756 18748
rect 23339 18717 23351 18720
rect 23293 18711 23351 18717
rect 22020 18680 22048 18711
rect 22204 18680 22232 18711
rect 23750 18708 23756 18720
rect 23808 18708 23814 18760
rect 24029 18751 24087 18757
rect 24029 18717 24041 18751
rect 24075 18748 24087 18751
rect 25130 18748 25136 18760
rect 24075 18720 25136 18748
rect 24075 18717 24087 18720
rect 24029 18711 24087 18717
rect 25130 18708 25136 18720
rect 25188 18708 25194 18760
rect 25501 18751 25559 18757
rect 25501 18717 25513 18751
rect 25547 18717 25559 18751
rect 25501 18711 25559 18717
rect 25593 18751 25651 18757
rect 25593 18717 25605 18751
rect 25639 18748 25651 18751
rect 25774 18748 25780 18760
rect 25639 18720 25780 18748
rect 25639 18717 25651 18720
rect 25593 18711 25651 18717
rect 23201 18683 23259 18689
rect 23201 18680 23213 18683
rect 22020 18652 22094 18680
rect 22204 18652 23213 18680
rect 22066 18612 22094 18652
rect 23201 18649 23213 18652
rect 23247 18649 23259 18683
rect 25516 18680 25544 18711
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18748 29055 18751
rect 29270 18748 29276 18760
rect 29043 18720 29276 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 29270 18708 29276 18720
rect 29328 18708 29334 18760
rect 30374 18748 30380 18760
rect 30335 18720 30380 18748
rect 30374 18708 30380 18720
rect 30432 18708 30438 18760
rect 31757 18751 31815 18757
rect 31757 18717 31769 18751
rect 31803 18717 31815 18751
rect 31757 18711 31815 18717
rect 32033 18751 32091 18757
rect 32033 18717 32045 18751
rect 32079 18748 32091 18751
rect 32122 18748 32128 18760
rect 32079 18720 32128 18748
rect 32079 18717 32091 18720
rect 32033 18711 32091 18717
rect 25682 18680 25688 18692
rect 25516 18652 25688 18680
rect 23201 18643 23259 18649
rect 25682 18640 25688 18652
rect 25740 18680 25746 18692
rect 26237 18683 26295 18689
rect 26237 18680 26249 18683
rect 25740 18652 26249 18680
rect 25740 18640 25746 18652
rect 26237 18649 26249 18652
rect 26283 18649 26295 18683
rect 26418 18680 26424 18692
rect 26379 18652 26424 18680
rect 26237 18643 26295 18649
rect 26418 18640 26424 18652
rect 26476 18640 26482 18692
rect 29086 18640 29092 18692
rect 29144 18680 29150 18692
rect 31772 18680 31800 18711
rect 32122 18708 32128 18720
rect 32180 18708 32186 18760
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32674 18748 32680 18760
rect 32272 18720 32680 18748
rect 32272 18708 32278 18720
rect 32674 18708 32680 18720
rect 32732 18708 32738 18760
rect 29144 18652 31800 18680
rect 29144 18640 29150 18652
rect 22278 18612 22284 18624
rect 22066 18584 22284 18612
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 23900 18584 24593 18612
rect 23900 18572 23906 18584
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 24581 18575 24639 18581
rect 25590 18572 25596 18624
rect 25648 18612 25654 18624
rect 25777 18615 25835 18621
rect 25777 18612 25789 18615
rect 25648 18584 25789 18612
rect 25648 18572 25654 18584
rect 25777 18581 25789 18584
rect 25823 18581 25835 18615
rect 31772 18612 31800 18652
rect 31941 18683 31999 18689
rect 31941 18649 31953 18683
rect 31987 18680 31999 18683
rect 32876 18680 32904 18779
rect 33226 18776 33232 18788
rect 33284 18776 33290 18828
rect 34514 18776 34520 18828
rect 34572 18816 34578 18828
rect 35802 18816 35808 18828
rect 34572 18788 35388 18816
rect 35763 18788 35808 18816
rect 34572 18776 34578 18788
rect 35360 18757 35388 18788
rect 35802 18776 35808 18788
rect 35860 18776 35866 18828
rect 36924 18760 36952 18856
rect 38654 18816 38660 18828
rect 37660 18788 38660 18816
rect 32953 18751 33011 18757
rect 32953 18717 32965 18751
rect 32999 18717 33011 18751
rect 32953 18711 33011 18717
rect 35161 18751 35219 18757
rect 35161 18717 35173 18751
rect 35207 18717 35219 18751
rect 35161 18711 35219 18717
rect 35345 18751 35403 18757
rect 35345 18717 35357 18751
rect 35391 18717 35403 18751
rect 35986 18748 35992 18760
rect 35947 18720 35992 18748
rect 35345 18711 35403 18717
rect 31987 18652 32904 18680
rect 31987 18649 31999 18652
rect 31941 18643 31999 18649
rect 32968 18612 32996 18711
rect 35176 18680 35204 18711
rect 35986 18708 35992 18720
rect 36044 18708 36050 18760
rect 36173 18751 36231 18757
rect 36173 18717 36185 18751
rect 36219 18748 36231 18751
rect 36722 18748 36728 18760
rect 36219 18720 36728 18748
rect 36219 18717 36231 18720
rect 36173 18711 36231 18717
rect 36722 18708 36728 18720
rect 36780 18708 36786 18760
rect 36906 18748 36912 18760
rect 36867 18720 36912 18748
rect 36906 18708 36912 18720
rect 36964 18708 36970 18760
rect 35618 18680 35624 18692
rect 35176 18652 35624 18680
rect 35618 18640 35624 18652
rect 35676 18640 35682 18692
rect 37660 18680 37688 18788
rect 38654 18776 38660 18788
rect 38712 18776 38718 18828
rect 38948 18816 38976 18856
rect 39022 18844 39028 18896
rect 39080 18884 39086 18896
rect 39117 18887 39175 18893
rect 39117 18884 39129 18887
rect 39080 18856 39129 18884
rect 39080 18844 39086 18856
rect 39117 18853 39129 18856
rect 39163 18853 39175 18887
rect 39117 18847 39175 18853
rect 45002 18844 45008 18896
rect 45060 18884 45066 18896
rect 45060 18856 51856 18884
rect 45060 18844 45066 18856
rect 39390 18816 39396 18828
rect 38948 18788 39396 18816
rect 39390 18776 39396 18788
rect 39448 18776 39454 18828
rect 40126 18816 40132 18828
rect 40087 18788 40132 18816
rect 40126 18776 40132 18788
rect 40184 18776 40190 18828
rect 40218 18776 40224 18828
rect 40276 18816 40282 18828
rect 40497 18819 40555 18825
rect 40497 18816 40509 18819
rect 40276 18788 40509 18816
rect 40276 18776 40282 18788
rect 40497 18785 40509 18788
rect 40543 18816 40555 18819
rect 41509 18819 41567 18825
rect 40543 18788 41460 18816
rect 40543 18785 40555 18788
rect 40497 18779 40555 18785
rect 38841 18751 38899 18757
rect 38841 18748 38853 18751
rect 38028 18720 38853 18748
rect 37826 18680 37832 18692
rect 36740 18652 37688 18680
rect 37787 18652 37832 18680
rect 36740 18624 36768 18652
rect 37826 18640 37832 18652
rect 37884 18640 37890 18692
rect 38028 18689 38056 18720
rect 38841 18717 38853 18720
rect 38887 18717 38899 18751
rect 38841 18711 38899 18717
rect 38979 18751 39037 18757
rect 38979 18717 38991 18751
rect 39025 18748 39037 18751
rect 39206 18748 39212 18760
rect 39025 18720 39212 18748
rect 39025 18717 39037 18720
rect 38979 18711 39037 18717
rect 38013 18683 38071 18689
rect 38013 18649 38025 18683
rect 38059 18649 38071 18683
rect 38856 18680 38884 18711
rect 39206 18708 39212 18720
rect 39264 18708 39270 18760
rect 39298 18708 39304 18760
rect 39356 18748 39362 18760
rect 40586 18748 40592 18760
rect 39356 18720 39401 18748
rect 40547 18720 40592 18748
rect 39356 18708 39362 18720
rect 40586 18708 40592 18720
rect 40644 18708 40650 18760
rect 41432 18757 41460 18788
rect 41509 18785 41521 18819
rect 41555 18785 41567 18819
rect 41782 18816 41788 18828
rect 41743 18788 41788 18816
rect 41509 18779 41567 18785
rect 41417 18751 41475 18757
rect 41417 18717 41429 18751
rect 41463 18717 41475 18751
rect 41417 18711 41475 18717
rect 39574 18680 39580 18692
rect 38856 18652 39580 18680
rect 38013 18643 38071 18649
rect 36630 18612 36636 18624
rect 31772 18584 36636 18612
rect 25777 18575 25835 18581
rect 36630 18572 36636 18584
rect 36688 18572 36694 18624
rect 36722 18572 36728 18624
rect 36780 18612 36786 18624
rect 36780 18584 36825 18612
rect 36780 18572 36786 18584
rect 37366 18572 37372 18624
rect 37424 18612 37430 18624
rect 38028 18612 38056 18643
rect 39574 18640 39580 18652
rect 39632 18640 39638 18692
rect 40604 18680 40632 18708
rect 41524 18680 41552 18779
rect 41782 18776 41788 18788
rect 41840 18776 41846 18828
rect 43441 18819 43499 18825
rect 43441 18785 43453 18819
rect 43487 18816 43499 18819
rect 45738 18816 45744 18828
rect 43487 18788 45744 18816
rect 43487 18785 43499 18788
rect 43441 18779 43499 18785
rect 45738 18776 45744 18788
rect 45796 18776 45802 18828
rect 46382 18776 46388 18828
rect 46440 18816 46446 18828
rect 49694 18816 49700 18828
rect 46440 18788 49700 18816
rect 46440 18776 46446 18788
rect 49694 18776 49700 18788
rect 49752 18776 49758 18828
rect 50525 18819 50583 18825
rect 50525 18785 50537 18819
rect 50571 18816 50583 18819
rect 50982 18816 50988 18828
rect 50571 18788 50988 18816
rect 50571 18785 50583 18788
rect 50525 18779 50583 18785
rect 50982 18776 50988 18788
rect 51040 18776 51046 18828
rect 51828 18816 51856 18856
rect 51902 18844 51908 18896
rect 51960 18884 51966 18896
rect 51960 18856 55812 18884
rect 51960 18844 51966 18856
rect 55784 18828 55812 18856
rect 52733 18819 52791 18825
rect 51828 18788 52684 18816
rect 43165 18751 43223 18757
rect 43165 18717 43177 18751
rect 43211 18748 43223 18751
rect 43254 18748 43260 18760
rect 43211 18720 43260 18748
rect 43211 18717 43223 18720
rect 43165 18711 43223 18717
rect 43254 18708 43260 18720
rect 43312 18708 43318 18760
rect 46661 18751 46719 18757
rect 46661 18717 46673 18751
rect 46707 18748 46719 18751
rect 46750 18748 46756 18760
rect 46707 18720 46756 18748
rect 46707 18717 46719 18720
rect 46661 18711 46719 18717
rect 46676 18680 46704 18711
rect 46750 18708 46756 18720
rect 46808 18708 46814 18760
rect 46934 18748 46940 18760
rect 46895 18720 46940 18748
rect 46934 18708 46940 18720
rect 46992 18748 46998 18760
rect 47397 18751 47455 18757
rect 47397 18748 47409 18751
rect 46992 18720 47409 18748
rect 46992 18708 46998 18720
rect 47397 18717 47409 18720
rect 47443 18717 47455 18751
rect 47578 18748 47584 18760
rect 47539 18720 47584 18748
rect 47397 18711 47455 18717
rect 47578 18708 47584 18720
rect 47636 18708 47642 18760
rect 50154 18708 50160 18760
rect 50212 18748 50218 18760
rect 50617 18751 50675 18757
rect 50617 18748 50629 18751
rect 50212 18720 50629 18748
rect 50212 18708 50218 18720
rect 50617 18717 50629 18720
rect 50663 18717 50675 18751
rect 50617 18711 50675 18717
rect 50706 18708 50712 18760
rect 50764 18748 50770 18760
rect 52089 18751 52147 18757
rect 50764 18720 50809 18748
rect 50764 18708 50770 18720
rect 52089 18717 52101 18751
rect 52135 18717 52147 18751
rect 52089 18711 52147 18717
rect 52365 18751 52423 18757
rect 52365 18717 52377 18751
rect 52411 18748 52423 18751
rect 52454 18748 52460 18760
rect 52411 18720 52460 18748
rect 52411 18717 52423 18720
rect 52365 18711 52423 18717
rect 40604 18652 41552 18680
rect 43272 18652 46704 18680
rect 46845 18683 46903 18689
rect 37424 18584 38056 18612
rect 37424 18572 37430 18584
rect 43162 18572 43168 18624
rect 43220 18612 43226 18624
rect 43272 18621 43300 18652
rect 46845 18649 46857 18683
rect 46891 18680 46903 18683
rect 47596 18680 47624 18708
rect 46891 18652 47624 18680
rect 52104 18680 52132 18711
rect 52454 18708 52460 18720
rect 52512 18708 52518 18760
rect 52656 18748 52684 18788
rect 52733 18785 52745 18819
rect 52779 18816 52791 18819
rect 52914 18816 52920 18828
rect 52779 18788 52920 18816
rect 52779 18785 52791 18788
rect 52733 18779 52791 18785
rect 52914 18776 52920 18788
rect 52972 18776 52978 18828
rect 55766 18816 55772 18828
rect 53576 18788 55076 18816
rect 55679 18788 55772 18816
rect 53576 18748 53604 18788
rect 52656 18720 53604 18748
rect 53653 18751 53711 18757
rect 53653 18717 53665 18751
rect 53699 18717 53711 18751
rect 53653 18711 53711 18717
rect 53668 18680 53696 18711
rect 54018 18708 54024 18760
rect 54076 18708 54082 18760
rect 52104 18652 53696 18680
rect 46891 18649 46903 18652
rect 46845 18643 46903 18649
rect 43257 18615 43315 18621
rect 43257 18612 43269 18615
rect 43220 18584 43269 18612
rect 43220 18572 43226 18584
rect 43257 18581 43269 18584
rect 43303 18581 43315 18615
rect 43257 18575 43315 18581
rect 43990 18572 43996 18624
rect 44048 18612 44054 18624
rect 44085 18615 44143 18621
rect 44085 18612 44097 18615
rect 44048 18584 44097 18612
rect 44048 18572 44054 18584
rect 44085 18581 44097 18584
rect 44131 18581 44143 18615
rect 44085 18575 44143 18581
rect 45281 18615 45339 18621
rect 45281 18581 45293 18615
rect 45327 18612 45339 18615
rect 45738 18612 45744 18624
rect 45327 18584 45744 18612
rect 45327 18581 45339 18584
rect 45281 18575 45339 18581
rect 45738 18572 45744 18584
rect 45796 18572 45802 18624
rect 45922 18612 45928 18624
rect 45883 18584 45928 18612
rect 45922 18572 45928 18584
rect 45980 18572 45986 18624
rect 47210 18572 47216 18624
rect 47268 18612 47274 18624
rect 48041 18615 48099 18621
rect 48041 18612 48053 18615
rect 47268 18584 48053 18612
rect 47268 18572 47274 18584
rect 48041 18581 48053 18584
rect 48087 18581 48099 18615
rect 48041 18575 48099 18581
rect 48685 18615 48743 18621
rect 48685 18581 48697 18615
rect 48731 18612 48743 18615
rect 49237 18615 49295 18621
rect 49237 18612 49249 18615
rect 48731 18584 49249 18612
rect 48731 18581 48743 18584
rect 48685 18575 48743 18581
rect 49237 18581 49249 18584
rect 49283 18612 49295 18615
rect 49789 18615 49847 18621
rect 49789 18612 49801 18615
rect 49283 18584 49801 18612
rect 49283 18581 49295 18584
rect 49237 18575 49295 18581
rect 49789 18581 49801 18584
rect 49835 18612 49847 18615
rect 50154 18612 50160 18624
rect 49835 18584 50160 18612
rect 49835 18581 49847 18584
rect 49789 18575 49847 18581
rect 50154 18572 50160 18584
rect 50212 18572 50218 18624
rect 53668 18612 53696 18652
rect 53926 18640 53932 18692
rect 53984 18680 53990 18692
rect 54389 18683 54447 18689
rect 54389 18680 54401 18683
rect 53984 18652 54401 18680
rect 53984 18640 53990 18652
rect 54389 18649 54401 18652
rect 54435 18649 54447 18683
rect 55048 18680 55076 18788
rect 55766 18776 55772 18788
rect 55824 18776 55830 18828
rect 55122 18708 55128 18760
rect 55180 18748 55186 18760
rect 55677 18751 55735 18757
rect 55677 18748 55689 18751
rect 55180 18720 55689 18748
rect 55180 18708 55186 18720
rect 55677 18717 55689 18720
rect 55723 18717 55735 18751
rect 55677 18711 55735 18717
rect 58069 18751 58127 18757
rect 58069 18717 58081 18751
rect 58115 18748 58127 18751
rect 58342 18748 58348 18760
rect 58115 18720 58348 18748
rect 58115 18717 58127 18720
rect 58069 18711 58127 18717
rect 58342 18708 58348 18720
rect 58400 18708 58406 18760
rect 55950 18680 55956 18692
rect 55048 18652 55956 18680
rect 54389 18643 54447 18649
rect 55950 18640 55956 18652
rect 56008 18680 56014 18692
rect 56597 18683 56655 18689
rect 56597 18680 56609 18683
rect 56008 18652 56609 18680
rect 56008 18640 56014 18652
rect 56597 18649 56609 18652
rect 56643 18649 56655 18683
rect 56597 18643 56655 18649
rect 55674 18612 55680 18624
rect 53668 18584 55680 18612
rect 55674 18572 55680 18584
rect 55732 18572 55738 18624
rect 56042 18572 56048 18624
rect 56100 18612 56106 18624
rect 56137 18615 56195 18621
rect 56137 18612 56149 18615
rect 56100 18584 56149 18612
rect 56100 18572 56106 18584
rect 56137 18581 56149 18584
rect 56183 18581 56195 18615
rect 57238 18612 57244 18624
rect 57199 18584 57244 18612
rect 56137 18575 56195 18581
rect 57238 18572 57244 18584
rect 57296 18572 57302 18624
rect 58250 18612 58256 18624
rect 58211 18584 58256 18612
rect 58250 18572 58256 18584
rect 58308 18572 58314 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 22094 18408 22100 18420
rect 22066 18368 22100 18408
rect 22152 18368 22158 18420
rect 23934 18368 23940 18420
rect 23992 18408 23998 18420
rect 24489 18411 24547 18417
rect 24489 18408 24501 18411
rect 23992 18380 24501 18408
rect 23992 18368 23998 18380
rect 24489 18377 24501 18380
rect 24535 18377 24547 18411
rect 24489 18371 24547 18377
rect 24673 18411 24731 18417
rect 24673 18377 24685 18411
rect 24719 18408 24731 18411
rect 25038 18408 25044 18420
rect 24719 18380 25044 18408
rect 24719 18377 24731 18380
rect 24673 18371 24731 18377
rect 25038 18368 25044 18380
rect 25096 18368 25102 18420
rect 25777 18411 25835 18417
rect 25777 18377 25789 18411
rect 25823 18408 25835 18411
rect 26234 18408 26240 18420
rect 25823 18380 26240 18408
rect 25823 18377 25835 18380
rect 25777 18371 25835 18377
rect 26234 18368 26240 18380
rect 26292 18368 26298 18420
rect 26326 18368 26332 18420
rect 26384 18408 26390 18420
rect 26605 18411 26663 18417
rect 26605 18408 26617 18411
rect 26384 18380 26617 18408
rect 26384 18368 26390 18380
rect 26605 18377 26617 18380
rect 26651 18377 26663 18411
rect 26605 18371 26663 18377
rect 27890 18368 27896 18420
rect 27948 18408 27954 18420
rect 28353 18411 28411 18417
rect 28353 18408 28365 18411
rect 27948 18380 28365 18408
rect 27948 18368 27954 18380
rect 28353 18377 28365 18380
rect 28399 18377 28411 18411
rect 30006 18408 30012 18420
rect 29967 18380 30012 18408
rect 28353 18371 28411 18377
rect 30006 18368 30012 18380
rect 30064 18368 30070 18420
rect 31110 18368 31116 18420
rect 31168 18408 31174 18420
rect 35250 18408 35256 18420
rect 31168 18380 35256 18408
rect 31168 18368 31174 18380
rect 35250 18368 35256 18380
rect 35308 18368 35314 18420
rect 35342 18368 35348 18420
rect 35400 18408 35406 18420
rect 35621 18411 35679 18417
rect 35621 18408 35633 18411
rect 35400 18380 35633 18408
rect 35400 18368 35406 18380
rect 35621 18377 35633 18380
rect 35667 18377 35679 18411
rect 35621 18371 35679 18377
rect 35805 18411 35863 18417
rect 35805 18377 35817 18411
rect 35851 18408 35863 18411
rect 36722 18408 36728 18420
rect 35851 18380 36728 18408
rect 35851 18377 35863 18380
rect 35805 18371 35863 18377
rect 36722 18368 36728 18380
rect 36780 18368 36786 18420
rect 38010 18368 38016 18420
rect 38068 18408 38074 18420
rect 38289 18411 38347 18417
rect 38289 18408 38301 18411
rect 38068 18380 38301 18408
rect 38068 18368 38074 18380
rect 38289 18377 38301 18380
rect 38335 18377 38347 18411
rect 38289 18371 38347 18377
rect 39761 18411 39819 18417
rect 39761 18377 39773 18411
rect 39807 18408 39819 18411
rect 40126 18408 40132 18420
rect 39807 18380 40132 18408
rect 39807 18377 39819 18380
rect 39761 18371 39819 18377
rect 40126 18368 40132 18380
rect 40184 18368 40190 18420
rect 41138 18368 41144 18420
rect 41196 18408 41202 18420
rect 41233 18411 41291 18417
rect 41233 18408 41245 18411
rect 41196 18380 41245 18408
rect 41196 18368 41202 18380
rect 41233 18377 41245 18380
rect 41279 18377 41291 18411
rect 41233 18371 41291 18377
rect 44085 18411 44143 18417
rect 44085 18377 44097 18411
rect 44131 18408 44143 18411
rect 44266 18408 44272 18420
rect 44131 18380 44272 18408
rect 44131 18377 44143 18380
rect 44085 18371 44143 18377
rect 44266 18368 44272 18380
rect 44324 18368 44330 18420
rect 52178 18408 52184 18420
rect 46216 18380 52184 18408
rect 22066 18340 22094 18368
rect 23842 18340 23848 18352
rect 22020 18312 22094 18340
rect 23506 18312 23848 18340
rect 1578 18272 1584 18284
rect 1539 18244 1584 18272
rect 1578 18232 1584 18244
rect 1636 18232 1642 18284
rect 22020 18281 22048 18312
rect 23842 18300 23848 18312
rect 23900 18300 23906 18352
rect 24854 18340 24860 18352
rect 24815 18312 24860 18340
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 25516 18312 26372 18340
rect 25516 18284 25544 18312
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 24762 18232 24768 18284
rect 24820 18272 24826 18284
rect 25041 18275 25099 18281
rect 24820 18244 24865 18272
rect 24820 18232 24826 18244
rect 25041 18241 25053 18275
rect 25087 18272 25099 18275
rect 25130 18272 25136 18284
rect 25087 18244 25136 18272
rect 25087 18241 25099 18244
rect 25041 18235 25099 18241
rect 22278 18204 22284 18216
rect 22191 18176 22284 18204
rect 22278 18164 22284 18176
rect 22336 18204 22342 18216
rect 23290 18204 23296 18216
rect 22336 18176 23296 18204
rect 22336 18164 22342 18176
rect 23290 18164 23296 18176
rect 23348 18164 23354 18216
rect 24029 18207 24087 18213
rect 24029 18173 24041 18207
rect 24075 18204 24087 18207
rect 25056 18204 25084 18235
rect 25130 18232 25136 18244
rect 25188 18232 25194 18284
rect 25498 18272 25504 18284
rect 25411 18244 25504 18272
rect 25498 18232 25504 18244
rect 25556 18232 25562 18284
rect 25590 18232 25596 18284
rect 25648 18272 25654 18284
rect 26234 18272 26240 18284
rect 25648 18244 25693 18272
rect 26195 18244 26240 18272
rect 25648 18232 25654 18244
rect 26234 18232 26240 18244
rect 26292 18232 26298 18284
rect 24075 18176 25084 18204
rect 24075 18173 24087 18176
rect 24029 18167 24087 18173
rect 25608 18136 25636 18232
rect 25777 18207 25835 18213
rect 25777 18173 25789 18207
rect 25823 18204 25835 18207
rect 26252 18204 26280 18232
rect 26344 18213 26372 18312
rect 26418 18300 26424 18352
rect 26476 18340 26482 18352
rect 27249 18343 27307 18349
rect 27249 18340 27261 18343
rect 26476 18312 27261 18340
rect 26476 18300 26482 18312
rect 27249 18309 27261 18312
rect 27295 18340 27307 18343
rect 37366 18340 37372 18352
rect 27295 18312 37372 18340
rect 27295 18309 27307 18312
rect 27249 18303 27307 18309
rect 37366 18300 37372 18312
rect 37424 18300 37430 18352
rect 37461 18343 37519 18349
rect 37461 18309 37473 18343
rect 37507 18340 37519 18343
rect 41782 18340 41788 18352
rect 37507 18312 38240 18340
rect 37507 18309 37519 18312
rect 37461 18303 37519 18309
rect 27154 18272 27160 18284
rect 27067 18244 27160 18272
rect 27154 18232 27160 18244
rect 27212 18272 27218 18284
rect 27985 18275 28043 18281
rect 27985 18272 27997 18275
rect 27212 18244 27997 18272
rect 27212 18232 27218 18244
rect 27985 18241 27997 18244
rect 28031 18241 28043 18275
rect 28166 18272 28172 18284
rect 28127 18244 28172 18272
rect 27985 18235 28043 18241
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 29546 18272 29552 18284
rect 29507 18244 29552 18272
rect 29546 18232 29552 18244
rect 29604 18232 29610 18284
rect 29825 18275 29883 18281
rect 29825 18241 29837 18275
rect 29871 18272 29883 18275
rect 29914 18272 29920 18284
rect 29871 18244 29920 18272
rect 29871 18241 29883 18244
rect 29825 18235 29883 18241
rect 29914 18232 29920 18244
rect 29972 18232 29978 18284
rect 30466 18272 30472 18284
rect 30427 18244 30472 18272
rect 30466 18232 30472 18244
rect 30524 18272 30530 18284
rect 31110 18272 31116 18284
rect 30524 18244 31116 18272
rect 30524 18232 30530 18244
rect 31110 18232 31116 18244
rect 31168 18232 31174 18284
rect 32766 18232 32772 18284
rect 32824 18272 32830 18284
rect 32861 18275 32919 18281
rect 32861 18272 32873 18275
rect 32824 18244 32873 18272
rect 32824 18232 32830 18244
rect 32861 18241 32873 18244
rect 32907 18241 32919 18275
rect 32861 18235 32919 18241
rect 32950 18232 32956 18284
rect 33008 18272 33014 18284
rect 33134 18272 33140 18284
rect 33008 18244 33053 18272
rect 33095 18244 33140 18272
rect 33008 18232 33014 18244
rect 33134 18232 33140 18244
rect 33192 18232 33198 18284
rect 35746 18275 35804 18281
rect 35746 18272 35758 18275
rect 33244 18244 35758 18272
rect 25823 18176 26280 18204
rect 26329 18207 26387 18213
rect 25823 18173 25835 18176
rect 25777 18167 25835 18173
rect 26329 18173 26341 18207
rect 26375 18204 26387 18207
rect 27246 18204 27252 18216
rect 26375 18176 27252 18204
rect 26375 18173 26387 18176
rect 26329 18167 26387 18173
rect 27246 18164 27252 18176
rect 27304 18164 27310 18216
rect 27890 18204 27896 18216
rect 27851 18176 27896 18204
rect 27890 18164 27896 18176
rect 27948 18164 27954 18216
rect 28074 18164 28080 18216
rect 28132 18204 28138 18216
rect 30561 18207 30619 18213
rect 28132 18176 28177 18204
rect 28132 18164 28138 18176
rect 30561 18173 30573 18207
rect 30607 18204 30619 18207
rect 31846 18204 31852 18216
rect 30607 18176 31852 18204
rect 30607 18173 30619 18176
rect 30561 18167 30619 18173
rect 31846 18164 31852 18176
rect 31904 18164 31910 18216
rect 32214 18164 32220 18216
rect 32272 18204 32278 18216
rect 33244 18204 33272 18244
rect 35746 18241 35758 18244
rect 35792 18241 35804 18275
rect 35746 18235 35804 18241
rect 36173 18275 36231 18281
rect 36173 18241 36185 18275
rect 36219 18272 36231 18275
rect 36538 18272 36544 18284
rect 36219 18244 36544 18272
rect 36219 18241 36231 18244
rect 36173 18235 36231 18241
rect 36538 18232 36544 18244
rect 36596 18232 36602 18284
rect 36630 18232 36636 18284
rect 36688 18272 36694 18284
rect 38212 18281 38240 18312
rect 41248 18312 41788 18340
rect 37737 18275 37795 18281
rect 37737 18272 37749 18275
rect 36688 18244 37749 18272
rect 36688 18232 36694 18244
rect 37737 18241 37749 18244
rect 37783 18241 37795 18275
rect 37737 18235 37795 18241
rect 38197 18275 38255 18281
rect 38197 18241 38209 18275
rect 38243 18241 38255 18275
rect 38378 18272 38384 18284
rect 38339 18244 38384 18272
rect 38197 18235 38255 18241
rect 38378 18232 38384 18244
rect 38436 18232 38442 18284
rect 39022 18232 39028 18284
rect 39080 18272 39086 18284
rect 39301 18275 39359 18281
rect 39301 18272 39313 18275
rect 39080 18244 39313 18272
rect 39080 18232 39086 18244
rect 39301 18241 39313 18244
rect 39347 18241 39359 18275
rect 39574 18272 39580 18284
rect 39535 18244 39580 18272
rect 39301 18235 39359 18241
rect 39574 18232 39580 18244
rect 39632 18232 39638 18284
rect 41248 18281 41276 18312
rect 41782 18300 41788 18312
rect 41840 18300 41846 18352
rect 41233 18275 41291 18281
rect 41233 18241 41245 18275
rect 41279 18241 41291 18275
rect 41233 18235 41291 18241
rect 41414 18232 41420 18284
rect 41472 18272 41478 18284
rect 42797 18275 42855 18281
rect 41472 18244 41517 18272
rect 41472 18232 41478 18244
rect 42797 18241 42809 18275
rect 42843 18272 42855 18275
rect 43349 18275 43407 18281
rect 43349 18272 43361 18275
rect 42843 18244 43361 18272
rect 42843 18241 42855 18244
rect 42797 18235 42855 18241
rect 43349 18241 43361 18244
rect 43395 18272 43407 18275
rect 43714 18272 43720 18284
rect 43395 18244 43720 18272
rect 43395 18241 43407 18244
rect 43349 18235 43407 18241
rect 43714 18232 43720 18244
rect 43772 18272 43778 18284
rect 43809 18275 43867 18281
rect 43809 18272 43821 18275
rect 43772 18244 43821 18272
rect 43772 18232 43778 18244
rect 43809 18241 43821 18244
rect 43855 18241 43867 18275
rect 43809 18235 43867 18241
rect 44450 18232 44456 18284
rect 44508 18272 44514 18284
rect 44729 18275 44787 18281
rect 44729 18272 44741 18275
rect 44508 18244 44741 18272
rect 44508 18232 44514 18244
rect 44729 18241 44741 18244
rect 44775 18241 44787 18275
rect 45646 18272 45652 18284
rect 45607 18244 45652 18272
rect 44729 18235 44787 18241
rect 45646 18232 45652 18244
rect 45704 18232 45710 18284
rect 46216 18281 46244 18380
rect 52178 18368 52184 18380
rect 52236 18368 52242 18420
rect 52822 18368 52828 18420
rect 52880 18408 52886 18420
rect 53377 18411 53435 18417
rect 53377 18408 53389 18411
rect 52880 18380 53389 18408
rect 52880 18368 52886 18380
rect 53377 18377 53389 18380
rect 53423 18377 53435 18411
rect 55122 18408 55128 18420
rect 55083 18380 55128 18408
rect 53377 18371 53435 18377
rect 55122 18368 55128 18380
rect 55180 18368 55186 18420
rect 46382 18340 46388 18352
rect 46343 18312 46388 18340
rect 46382 18300 46388 18312
rect 46440 18300 46446 18352
rect 50706 18340 50712 18352
rect 46860 18312 50712 18340
rect 45833 18275 45891 18281
rect 45833 18241 45845 18275
rect 45879 18241 45891 18275
rect 45833 18235 45891 18241
rect 45925 18275 45983 18281
rect 45925 18241 45937 18275
rect 45971 18272 45983 18275
rect 46201 18275 46259 18281
rect 45971 18244 46152 18272
rect 45971 18241 45983 18244
rect 45925 18235 45983 18241
rect 32272 18176 33272 18204
rect 36265 18207 36323 18213
rect 32272 18164 32278 18176
rect 36265 18173 36277 18207
rect 36311 18204 36323 18207
rect 36722 18204 36728 18216
rect 36311 18176 36728 18204
rect 36311 18173 36323 18176
rect 36265 18167 36323 18173
rect 36722 18164 36728 18176
rect 36780 18164 36786 18216
rect 37458 18204 37464 18216
rect 37419 18176 37464 18204
rect 37458 18164 37464 18176
rect 37516 18164 37522 18216
rect 39206 18164 39212 18216
rect 39264 18204 39270 18216
rect 39393 18207 39451 18213
rect 39393 18204 39405 18207
rect 39264 18176 39405 18204
rect 39264 18164 39270 18176
rect 39393 18173 39405 18176
rect 39439 18173 39451 18207
rect 39393 18167 39451 18173
rect 44085 18207 44143 18213
rect 44085 18173 44097 18207
rect 44131 18204 44143 18207
rect 44542 18204 44548 18216
rect 44131 18176 44548 18204
rect 44131 18173 44143 18176
rect 44085 18167 44143 18173
rect 44542 18164 44548 18176
rect 44600 18164 44606 18216
rect 44637 18207 44695 18213
rect 44637 18173 44649 18207
rect 44683 18173 44695 18207
rect 44637 18167 44695 18173
rect 29638 18136 29644 18148
rect 25608 18108 26280 18136
rect 29599 18108 29644 18136
rect 1762 18068 1768 18080
rect 1723 18040 1768 18068
rect 1762 18028 1768 18040
rect 1820 18028 1826 18080
rect 26252 18077 26280 18108
rect 29638 18096 29644 18108
rect 29696 18096 29702 18148
rect 29733 18139 29791 18145
rect 29733 18105 29745 18139
rect 29779 18136 29791 18139
rect 29822 18136 29828 18148
rect 29779 18108 29828 18136
rect 29779 18105 29791 18108
rect 29733 18099 29791 18105
rect 29822 18096 29828 18108
rect 29880 18096 29886 18148
rect 33137 18139 33195 18145
rect 33137 18105 33149 18139
rect 33183 18136 33195 18139
rect 44652 18136 44680 18167
rect 44818 18164 44824 18216
rect 44876 18204 44882 18216
rect 45848 18204 45876 18235
rect 44876 18176 45876 18204
rect 46017 18207 46075 18213
rect 44876 18164 44882 18176
rect 46017 18173 46029 18207
rect 46063 18173 46075 18207
rect 46124 18204 46152 18244
rect 46201 18241 46213 18275
rect 46247 18241 46259 18275
rect 46201 18235 46259 18241
rect 46860 18213 46888 18312
rect 50706 18300 50712 18312
rect 50764 18300 50770 18352
rect 53742 18340 53748 18352
rect 53703 18312 53748 18340
rect 53742 18300 53748 18312
rect 53800 18300 53806 18352
rect 55674 18340 55680 18352
rect 55635 18312 55680 18340
rect 55674 18300 55680 18312
rect 55732 18300 55738 18352
rect 48317 18275 48375 18281
rect 48317 18241 48329 18275
rect 48363 18241 48375 18275
rect 48498 18272 48504 18284
rect 48459 18244 48504 18272
rect 48317 18235 48375 18241
rect 46845 18207 46903 18213
rect 46845 18204 46857 18207
rect 46124 18176 46857 18204
rect 46017 18167 46075 18173
rect 46845 18173 46857 18176
rect 46891 18173 46903 18207
rect 48332 18204 48360 18235
rect 48498 18232 48504 18244
rect 48556 18232 48562 18284
rect 48958 18272 48964 18284
rect 48919 18244 48964 18272
rect 48958 18232 48964 18244
rect 49016 18232 49022 18284
rect 49145 18275 49203 18281
rect 49145 18241 49157 18275
rect 49191 18272 49203 18275
rect 50154 18272 50160 18284
rect 49191 18244 50160 18272
rect 49191 18241 49203 18244
rect 49145 18235 49203 18241
rect 50154 18232 50160 18244
rect 50212 18232 50218 18284
rect 50341 18275 50399 18281
rect 50341 18241 50353 18275
rect 50387 18272 50399 18275
rect 51902 18272 51908 18284
rect 50387 18244 51908 18272
rect 50387 18241 50399 18244
rect 50341 18235 50399 18241
rect 51902 18232 51908 18244
rect 51960 18232 51966 18284
rect 53561 18275 53619 18281
rect 53561 18241 53573 18275
rect 53607 18241 53619 18275
rect 53561 18235 53619 18241
rect 49053 18207 49111 18213
rect 49053 18204 49065 18207
rect 48332 18176 49065 18204
rect 46845 18167 46903 18173
rect 49053 18173 49065 18176
rect 49099 18204 49111 18207
rect 51166 18204 51172 18216
rect 49099 18176 51172 18204
rect 49099 18173 49111 18176
rect 49053 18167 49111 18173
rect 45002 18136 45008 18148
rect 33183 18108 38654 18136
rect 44652 18108 45008 18136
rect 33183 18105 33195 18108
rect 33137 18099 33195 18105
rect 26237 18071 26295 18077
rect 26237 18037 26249 18071
rect 26283 18037 26295 18071
rect 26237 18031 26295 18037
rect 27522 18028 27528 18080
rect 27580 18068 27586 18080
rect 28258 18068 28264 18080
rect 27580 18040 28264 18068
rect 27580 18028 27586 18040
rect 28258 18028 28264 18040
rect 28316 18028 28322 18080
rect 28534 18028 28540 18080
rect 28592 18068 28598 18080
rect 28902 18068 28908 18080
rect 28592 18040 28908 18068
rect 28592 18028 28598 18040
rect 28902 18028 28908 18040
rect 28960 18028 28966 18080
rect 35250 18028 35256 18080
rect 35308 18068 35314 18080
rect 36817 18071 36875 18077
rect 36817 18068 36829 18071
rect 35308 18040 36829 18068
rect 35308 18028 35314 18040
rect 36817 18037 36829 18040
rect 36863 18068 36875 18071
rect 36906 18068 36912 18080
rect 36863 18040 36912 18068
rect 36863 18037 36875 18040
rect 36817 18031 36875 18037
rect 36906 18028 36912 18040
rect 36964 18028 36970 18080
rect 37366 18028 37372 18080
rect 37424 18068 37430 18080
rect 37645 18071 37703 18077
rect 37645 18068 37657 18071
rect 37424 18040 37657 18068
rect 37424 18028 37430 18040
rect 37645 18037 37657 18040
rect 37691 18037 37703 18071
rect 38626 18068 38654 18108
rect 45002 18096 45008 18108
rect 45060 18096 45066 18148
rect 45097 18139 45155 18145
rect 45097 18105 45109 18139
rect 45143 18136 45155 18139
rect 46032 18136 46060 18167
rect 51166 18164 51172 18176
rect 51224 18164 51230 18216
rect 51442 18164 51448 18216
rect 51500 18204 51506 18216
rect 53576 18204 53604 18235
rect 53650 18232 53656 18284
rect 53708 18272 53714 18284
rect 53708 18244 53753 18272
rect 53708 18232 53714 18244
rect 53926 18232 53932 18284
rect 53984 18272 53990 18284
rect 55033 18275 55091 18281
rect 53984 18244 54029 18272
rect 53984 18232 53990 18244
rect 55033 18241 55045 18275
rect 55079 18241 55091 18275
rect 55766 18272 55772 18284
rect 55727 18244 55772 18272
rect 55033 18235 55091 18241
rect 55048 18204 55076 18235
rect 55766 18232 55772 18244
rect 55824 18232 55830 18284
rect 55950 18272 55956 18284
rect 55911 18244 55956 18272
rect 55950 18232 55956 18244
rect 56008 18272 56014 18284
rect 57057 18275 57115 18281
rect 57057 18272 57069 18275
rect 56008 18244 57069 18272
rect 56008 18232 56014 18244
rect 57057 18241 57069 18244
rect 57103 18272 57115 18275
rect 57790 18272 57796 18284
rect 57103 18244 57796 18272
rect 57103 18241 57115 18244
rect 57057 18235 57115 18241
rect 57790 18232 57796 18244
rect 57848 18272 57854 18284
rect 58069 18275 58127 18281
rect 58069 18272 58081 18275
rect 57848 18244 58081 18272
rect 57848 18232 57854 18244
rect 58069 18241 58081 18244
rect 58115 18241 58127 18275
rect 58069 18235 58127 18241
rect 51500 18176 55076 18204
rect 51500 18164 51506 18176
rect 45143 18108 46060 18136
rect 45143 18105 45155 18108
rect 45097 18099 45155 18105
rect 47578 18096 47584 18148
rect 47636 18136 47642 18148
rect 48317 18139 48375 18145
rect 48317 18136 48329 18139
rect 47636 18108 48329 18136
rect 47636 18096 47642 18108
rect 48317 18105 48329 18108
rect 48363 18105 48375 18139
rect 48317 18099 48375 18105
rect 49510 18096 49516 18148
rect 49568 18136 49574 18148
rect 49568 18108 50108 18136
rect 49568 18096 49574 18108
rect 39298 18068 39304 18080
rect 38626 18040 39304 18068
rect 37645 18031 37703 18037
rect 39298 18028 39304 18040
rect 39356 18028 39362 18080
rect 43898 18068 43904 18080
rect 43859 18040 43904 18068
rect 43898 18028 43904 18040
rect 43956 18028 43962 18080
rect 48041 18071 48099 18077
rect 48041 18037 48053 18071
rect 48087 18068 48099 18071
rect 48406 18068 48412 18080
rect 48087 18040 48412 18068
rect 48087 18037 48099 18040
rect 48041 18031 48099 18037
rect 48406 18028 48412 18040
rect 48464 18028 48470 18080
rect 49786 18028 49792 18080
rect 49844 18068 49850 18080
rect 49973 18071 50031 18077
rect 49973 18068 49985 18071
rect 49844 18040 49985 18068
rect 49844 18028 49850 18040
rect 49973 18037 49985 18040
rect 50019 18037 50031 18071
rect 50080 18068 50108 18108
rect 50154 18096 50160 18148
rect 50212 18136 50218 18148
rect 50890 18136 50896 18148
rect 50212 18108 50896 18136
rect 50212 18096 50218 18108
rect 50890 18096 50896 18108
rect 50948 18096 50954 18148
rect 54202 18096 54208 18148
rect 54260 18136 54266 18148
rect 56505 18139 56563 18145
rect 56505 18136 56517 18139
rect 54260 18108 56517 18136
rect 54260 18096 54266 18108
rect 56505 18105 56517 18108
rect 56551 18136 56563 18139
rect 57422 18136 57428 18148
rect 56551 18108 57428 18136
rect 56551 18105 56563 18108
rect 56505 18099 56563 18105
rect 57422 18096 57428 18108
rect 57480 18096 57486 18148
rect 51445 18071 51503 18077
rect 51445 18068 51457 18071
rect 50080 18040 51457 18068
rect 49973 18031 50031 18037
rect 51445 18037 51457 18040
rect 51491 18037 51503 18071
rect 51902 18068 51908 18080
rect 51863 18040 51908 18068
rect 51445 18031 51503 18037
rect 51902 18028 51908 18040
rect 51960 18028 51966 18080
rect 52362 18028 52368 18080
rect 52420 18068 52426 18080
rect 54389 18071 54447 18077
rect 54389 18068 54401 18071
rect 52420 18040 54401 18068
rect 52420 18028 52426 18040
rect 54389 18037 54401 18040
rect 54435 18068 54447 18071
rect 54754 18068 54760 18080
rect 54435 18040 54760 18068
rect 54435 18037 54447 18040
rect 54389 18031 54447 18037
rect 54754 18028 54760 18040
rect 54812 18028 54818 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 23290 17864 23296 17876
rect 23251 17836 23296 17864
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24581 17867 24639 17873
rect 24581 17864 24593 17867
rect 24084 17836 24593 17864
rect 24084 17824 24090 17836
rect 24581 17833 24593 17836
rect 24627 17833 24639 17867
rect 24581 17827 24639 17833
rect 24946 17824 24952 17876
rect 25004 17864 25010 17876
rect 25774 17864 25780 17876
rect 25004 17836 25780 17864
rect 25004 17824 25010 17836
rect 25774 17824 25780 17836
rect 25832 17864 25838 17876
rect 26329 17867 26387 17873
rect 26329 17864 26341 17867
rect 25832 17836 26341 17864
rect 25832 17824 25838 17836
rect 26329 17833 26341 17836
rect 26375 17833 26387 17867
rect 26329 17827 26387 17833
rect 27522 17824 27528 17876
rect 27580 17864 27586 17876
rect 27580 17836 27752 17864
rect 27580 17824 27586 17836
rect 1578 17796 1584 17808
rect 1539 17768 1584 17796
rect 1578 17756 1584 17768
rect 1636 17756 1642 17808
rect 23937 17799 23995 17805
rect 23937 17765 23949 17799
rect 23983 17796 23995 17799
rect 27246 17796 27252 17808
rect 23983 17768 24900 17796
rect 27159 17768 27252 17796
rect 23983 17765 23995 17768
rect 23937 17759 23995 17765
rect 24872 17740 24900 17768
rect 27246 17756 27252 17768
rect 27304 17796 27310 17808
rect 27724 17796 27752 17836
rect 27798 17824 27804 17876
rect 27856 17864 27862 17876
rect 28077 17867 28135 17873
rect 28077 17864 28089 17867
rect 27856 17836 28089 17864
rect 27856 17824 27862 17836
rect 28077 17833 28089 17836
rect 28123 17833 28135 17867
rect 28997 17867 29055 17873
rect 28997 17864 29009 17867
rect 28077 17827 28135 17833
rect 28184 17836 29009 17864
rect 28184 17796 28212 17836
rect 28997 17833 29009 17836
rect 29043 17864 29055 17867
rect 33226 17864 33232 17876
rect 29043 17836 33232 17864
rect 29043 17833 29055 17836
rect 28997 17827 29055 17833
rect 33226 17824 33232 17836
rect 33284 17824 33290 17876
rect 33778 17864 33784 17876
rect 33739 17836 33784 17864
rect 33778 17824 33784 17836
rect 33836 17824 33842 17876
rect 35253 17867 35311 17873
rect 35253 17833 35265 17867
rect 35299 17864 35311 17867
rect 35434 17864 35440 17876
rect 35299 17836 35440 17864
rect 35299 17833 35311 17836
rect 35253 17827 35311 17833
rect 35434 17824 35440 17836
rect 35492 17824 35498 17876
rect 36446 17824 36452 17876
rect 36504 17864 36510 17876
rect 36817 17867 36875 17873
rect 36817 17864 36829 17867
rect 36504 17836 36829 17864
rect 36504 17824 36510 17836
rect 36817 17833 36829 17836
rect 36863 17833 36875 17867
rect 38746 17864 38752 17876
rect 36817 17827 36875 17833
rect 37844 17836 38752 17864
rect 27304 17768 27660 17796
rect 27724 17768 28212 17796
rect 31297 17799 31355 17805
rect 27304 17756 27310 17768
rect 24026 17728 24032 17740
rect 23987 17700 24032 17728
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 24762 17728 24768 17740
rect 24723 17700 24768 17728
rect 24762 17688 24768 17700
rect 24820 17688 24826 17740
rect 24854 17688 24860 17740
rect 24912 17728 24918 17740
rect 24912 17700 24957 17728
rect 24912 17688 24918 17700
rect 23750 17660 23756 17672
rect 23711 17632 23756 17660
rect 23750 17620 23756 17632
rect 23808 17620 23814 17672
rect 23845 17663 23903 17669
rect 23845 17629 23857 17663
rect 23891 17660 23903 17663
rect 24949 17663 25007 17669
rect 23891 17632 24900 17660
rect 23891 17629 23903 17632
rect 23845 17623 23903 17629
rect 24872 17524 24900 17632
rect 24949 17629 24961 17663
rect 24995 17629 25007 17663
rect 24949 17623 25007 17629
rect 24964 17592 24992 17623
rect 25038 17620 25044 17672
rect 25096 17660 25102 17672
rect 26694 17660 26700 17672
rect 25096 17632 25141 17660
rect 26436 17632 26700 17660
rect 25096 17620 25102 17632
rect 25130 17592 25136 17604
rect 24964 17564 25136 17592
rect 25130 17552 25136 17564
rect 25188 17552 25194 17604
rect 25682 17592 25688 17604
rect 25240 17564 25688 17592
rect 25240 17524 25268 17564
rect 25682 17552 25688 17564
rect 25740 17592 25746 17604
rect 26145 17595 26203 17601
rect 26145 17592 26157 17595
rect 25740 17564 26157 17592
rect 25740 17552 25746 17564
rect 26145 17561 26157 17564
rect 26191 17561 26203 17595
rect 26145 17555 26203 17561
rect 26234 17552 26240 17604
rect 26292 17592 26298 17604
rect 26350 17595 26408 17601
rect 26350 17592 26362 17595
rect 26292 17564 26362 17592
rect 26292 17552 26298 17564
rect 26350 17561 26362 17564
rect 26396 17592 26408 17595
rect 26436 17592 26464 17632
rect 26694 17620 26700 17632
rect 26752 17620 26758 17672
rect 27264 17669 27292 17756
rect 27522 17728 27528 17740
rect 27483 17700 27528 17728
rect 27522 17688 27528 17700
rect 27580 17688 27586 17740
rect 27632 17728 27660 17768
rect 31297 17765 31309 17799
rect 31343 17796 31355 17799
rect 31386 17796 31392 17808
rect 31343 17768 31392 17796
rect 31343 17765 31355 17768
rect 31297 17759 31355 17765
rect 31386 17756 31392 17768
rect 31444 17756 31450 17808
rect 34514 17796 34520 17808
rect 33612 17768 34520 17796
rect 29086 17728 29092 17740
rect 27632 17700 29092 17728
rect 29086 17688 29092 17700
rect 29144 17688 29150 17740
rect 31021 17731 31079 17737
rect 31021 17697 31033 17731
rect 31067 17728 31079 17731
rect 31202 17728 31208 17740
rect 31067 17700 31208 17728
rect 31067 17697 31079 17700
rect 31021 17691 31079 17697
rect 31202 17688 31208 17700
rect 31260 17688 31266 17740
rect 32306 17688 32312 17740
rect 32364 17728 32370 17740
rect 33612 17728 33640 17768
rect 34514 17756 34520 17768
rect 34572 17756 34578 17808
rect 32364 17700 33640 17728
rect 32364 17688 32370 17700
rect 27249 17663 27307 17669
rect 27249 17629 27261 17663
rect 27295 17629 27307 17663
rect 27249 17623 27307 17629
rect 27341 17663 27399 17669
rect 27341 17629 27353 17663
rect 27387 17629 27399 17663
rect 27982 17660 27988 17672
rect 27943 17632 27988 17660
rect 27341 17623 27399 17629
rect 27356 17592 27384 17623
rect 27982 17620 27988 17632
rect 28040 17620 28046 17672
rect 28077 17663 28135 17669
rect 28077 17629 28089 17663
rect 28123 17660 28135 17663
rect 28166 17660 28172 17672
rect 28123 17632 28172 17660
rect 28123 17629 28135 17632
rect 28077 17623 28135 17629
rect 28166 17620 28172 17632
rect 28224 17620 28230 17672
rect 28258 17620 28264 17672
rect 28316 17660 28322 17672
rect 28353 17663 28411 17669
rect 28353 17660 28365 17663
rect 28316 17632 28365 17660
rect 28316 17620 28322 17632
rect 28353 17629 28365 17632
rect 28399 17629 28411 17663
rect 28353 17623 28411 17629
rect 29181 17663 29239 17669
rect 29181 17629 29193 17663
rect 29227 17629 29239 17663
rect 30926 17660 30932 17672
rect 30887 17632 30932 17660
rect 29181 17623 29239 17629
rect 29196 17592 29224 17623
rect 30926 17620 30932 17632
rect 30984 17620 30990 17672
rect 32398 17660 32404 17672
rect 32359 17632 32404 17660
rect 32398 17620 32404 17632
rect 32456 17620 32462 17672
rect 32585 17663 32643 17669
rect 32585 17629 32597 17663
rect 32631 17660 32643 17663
rect 32674 17660 32680 17672
rect 32631 17632 32680 17660
rect 32631 17629 32643 17632
rect 32585 17623 32643 17629
rect 32674 17620 32680 17632
rect 32732 17620 32738 17672
rect 32769 17663 32827 17669
rect 32769 17629 32781 17663
rect 32815 17629 32827 17663
rect 32769 17623 32827 17629
rect 33045 17663 33103 17669
rect 33045 17629 33057 17663
rect 33091 17629 33103 17663
rect 33045 17623 33103 17629
rect 33137 17663 33195 17669
rect 33137 17629 33149 17663
rect 33183 17660 33195 17663
rect 33226 17660 33232 17672
rect 33183 17632 33232 17660
rect 33183 17629 33195 17632
rect 33137 17623 33195 17629
rect 32122 17592 32128 17604
rect 26396 17564 26464 17592
rect 26528 17564 32128 17592
rect 26396 17561 26408 17564
rect 26350 17555 26408 17561
rect 25590 17524 25596 17536
rect 24872 17496 25268 17524
rect 25551 17496 25596 17524
rect 25590 17484 25596 17496
rect 25648 17484 25654 17536
rect 26528 17533 26556 17564
rect 32122 17552 32128 17564
rect 32180 17592 32186 17604
rect 32784 17592 32812 17623
rect 32180 17564 32812 17592
rect 33060 17592 33088 17623
rect 33226 17620 33232 17632
rect 33284 17620 33290 17672
rect 33612 17669 33640 17700
rect 33873 17731 33931 17737
rect 33873 17697 33885 17731
rect 33919 17728 33931 17731
rect 34054 17728 34060 17740
rect 33919 17700 34060 17728
rect 33919 17697 33931 17700
rect 33873 17691 33931 17697
rect 34054 17688 34060 17700
rect 34112 17728 34118 17740
rect 34885 17731 34943 17737
rect 34885 17728 34897 17731
rect 34112 17700 34897 17728
rect 34112 17688 34118 17700
rect 34885 17697 34897 17700
rect 34931 17697 34943 17731
rect 34885 17691 34943 17697
rect 37093 17731 37151 17737
rect 37093 17697 37105 17731
rect 37139 17728 37151 17731
rect 37734 17728 37740 17740
rect 37139 17700 37740 17728
rect 37139 17697 37151 17700
rect 37093 17691 37151 17697
rect 37734 17688 37740 17700
rect 37792 17688 37798 17740
rect 33597 17663 33655 17669
rect 33597 17629 33609 17663
rect 33643 17629 33655 17663
rect 33597 17623 33655 17629
rect 33686 17620 33692 17672
rect 33744 17660 33750 17672
rect 33744 17632 33789 17660
rect 33744 17620 33750 17632
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 35069 17663 35127 17669
rect 35069 17660 35081 17663
rect 34572 17632 35081 17660
rect 34572 17620 34578 17632
rect 35069 17629 35081 17632
rect 35115 17629 35127 17663
rect 35069 17623 35127 17629
rect 36630 17620 36636 17672
rect 36688 17660 36694 17672
rect 37001 17663 37059 17669
rect 37001 17660 37013 17663
rect 36688 17632 37013 17660
rect 36688 17620 36694 17632
rect 37001 17629 37013 17632
rect 37047 17629 37059 17663
rect 37182 17660 37188 17672
rect 37143 17632 37188 17660
rect 37001 17623 37059 17629
rect 37182 17620 37188 17632
rect 37240 17620 37246 17672
rect 37274 17620 37280 17672
rect 37332 17660 37338 17672
rect 37332 17632 37377 17660
rect 37332 17620 37338 17632
rect 37458 17620 37464 17672
rect 37516 17660 37522 17672
rect 37516 17632 37561 17660
rect 37516 17620 37522 17632
rect 37844 17592 37872 17836
rect 38746 17824 38752 17836
rect 38804 17864 38810 17876
rect 39025 17867 39083 17873
rect 39025 17864 39037 17867
rect 38804 17836 39037 17864
rect 38804 17824 38810 17836
rect 39025 17833 39037 17836
rect 39071 17833 39083 17867
rect 39206 17864 39212 17876
rect 39167 17836 39212 17864
rect 39025 17827 39083 17833
rect 39206 17824 39212 17836
rect 39264 17824 39270 17876
rect 44542 17824 44548 17876
rect 44600 17864 44606 17876
rect 45189 17867 45247 17873
rect 45189 17864 45201 17867
rect 44600 17836 45201 17864
rect 44600 17824 44606 17836
rect 45189 17833 45201 17836
rect 45235 17833 45247 17867
rect 45189 17827 45247 17833
rect 46014 17824 46020 17876
rect 46072 17864 46078 17876
rect 46072 17836 47072 17864
rect 46072 17824 46078 17836
rect 43901 17799 43959 17805
rect 43901 17765 43913 17799
rect 43947 17796 43959 17799
rect 44818 17796 44824 17808
rect 43947 17768 44824 17796
rect 43947 17765 43959 17768
rect 43901 17759 43959 17765
rect 44818 17756 44824 17768
rect 44876 17756 44882 17808
rect 46106 17756 46112 17808
rect 46164 17796 46170 17808
rect 47044 17796 47072 17836
rect 47486 17824 47492 17876
rect 47544 17864 47550 17876
rect 48409 17867 48467 17873
rect 48409 17864 48421 17867
rect 47544 17836 48421 17864
rect 47544 17824 47550 17836
rect 48409 17833 48421 17836
rect 48455 17833 48467 17867
rect 48409 17827 48467 17833
rect 47581 17799 47639 17805
rect 47581 17796 47593 17799
rect 46164 17768 46914 17796
rect 47044 17768 47593 17796
rect 46164 17756 46170 17768
rect 43533 17731 43591 17737
rect 43533 17697 43545 17731
rect 43579 17728 43591 17731
rect 44453 17731 44511 17737
rect 44453 17728 44465 17731
rect 43579 17700 44465 17728
rect 43579 17697 43591 17700
rect 43533 17691 43591 17697
rect 44453 17697 44465 17700
rect 44499 17728 44511 17731
rect 46886 17728 46914 17768
rect 47581 17765 47593 17768
rect 47627 17796 47639 17799
rect 47762 17796 47768 17808
rect 47627 17768 47768 17796
rect 47627 17765 47639 17768
rect 47581 17759 47639 17765
rect 47762 17756 47768 17768
rect 47820 17756 47826 17808
rect 48424 17796 48452 17827
rect 48498 17824 48504 17876
rect 48556 17864 48562 17876
rect 48593 17867 48651 17873
rect 48593 17864 48605 17867
rect 48556 17836 48605 17864
rect 48556 17824 48562 17836
rect 48593 17833 48605 17836
rect 48639 17833 48651 17867
rect 50982 17864 50988 17876
rect 50943 17836 50988 17864
rect 48593 17827 48651 17833
rect 50982 17824 50988 17836
rect 51040 17824 51046 17876
rect 51718 17824 51724 17876
rect 51776 17864 51782 17876
rect 51813 17867 51871 17873
rect 51813 17864 51825 17867
rect 51776 17836 51825 17864
rect 51776 17824 51782 17836
rect 51813 17833 51825 17836
rect 51859 17833 51871 17867
rect 51813 17827 51871 17833
rect 53098 17824 53104 17876
rect 53156 17864 53162 17876
rect 53193 17867 53251 17873
rect 53193 17864 53205 17867
rect 53156 17836 53205 17864
rect 53156 17824 53162 17836
rect 53193 17833 53205 17836
rect 53239 17833 53251 17867
rect 53193 17827 53251 17833
rect 53466 17824 53472 17876
rect 53524 17864 53530 17876
rect 53837 17867 53895 17873
rect 53837 17864 53849 17867
rect 53524 17836 53849 17864
rect 53524 17824 53530 17836
rect 53837 17833 53849 17836
rect 53883 17833 53895 17867
rect 53837 17827 53895 17833
rect 54205 17867 54263 17873
rect 54205 17833 54217 17867
rect 54251 17864 54263 17867
rect 54478 17864 54484 17876
rect 54251 17836 54484 17864
rect 54251 17833 54263 17836
rect 54205 17827 54263 17833
rect 54478 17824 54484 17836
rect 54536 17824 54542 17876
rect 55493 17867 55551 17873
rect 55493 17833 55505 17867
rect 55539 17864 55551 17867
rect 55582 17864 55588 17876
rect 55539 17836 55588 17864
rect 55539 17833 55551 17836
rect 55493 17827 55551 17833
rect 55582 17824 55588 17836
rect 55640 17824 55646 17876
rect 57790 17864 57796 17876
rect 57751 17836 57796 17864
rect 57790 17824 57796 17836
rect 57848 17824 57854 17876
rect 48958 17796 48964 17808
rect 48424 17768 48964 17796
rect 48958 17756 48964 17768
rect 49016 17756 49022 17808
rect 49605 17799 49663 17805
rect 49605 17765 49617 17799
rect 49651 17796 49663 17799
rect 52089 17799 52147 17805
rect 52089 17796 52101 17799
rect 49651 17768 50752 17796
rect 49651 17765 49663 17768
rect 49605 17759 49663 17765
rect 49786 17728 49792 17740
rect 44499 17700 46612 17728
rect 46886 17700 49648 17728
rect 49747 17700 49792 17728
rect 44499 17697 44511 17700
rect 44453 17691 44511 17697
rect 37921 17663 37979 17669
rect 37921 17629 37933 17663
rect 37967 17629 37979 17663
rect 37921 17623 37979 17629
rect 43257 17663 43315 17669
rect 43257 17629 43269 17663
rect 43303 17629 43315 17663
rect 43438 17660 43444 17672
rect 43399 17632 43444 17660
rect 43257 17623 43315 17629
rect 33060 17564 37872 17592
rect 32180 17552 32186 17564
rect 26513 17527 26571 17533
rect 26513 17493 26525 17527
rect 26559 17493 26571 17527
rect 26513 17487 26571 17493
rect 27525 17527 27583 17533
rect 27525 17493 27537 17527
rect 27571 17524 27583 17527
rect 28074 17524 28080 17536
rect 27571 17496 28080 17524
rect 27571 17493 27583 17496
rect 27525 17487 27583 17493
rect 28074 17484 28080 17496
rect 28132 17524 28138 17536
rect 28169 17527 28227 17533
rect 28169 17524 28181 17527
rect 28132 17496 28181 17524
rect 28132 17484 28138 17496
rect 28169 17493 28181 17496
rect 28215 17493 28227 17527
rect 28169 17487 28227 17493
rect 28258 17484 28264 17536
rect 28316 17524 28322 17536
rect 28813 17527 28871 17533
rect 28813 17524 28825 17527
rect 28316 17496 28825 17524
rect 28316 17484 28322 17496
rect 28813 17493 28825 17496
rect 28859 17493 28871 17527
rect 28813 17487 28871 17493
rect 36630 17484 36636 17536
rect 36688 17524 36694 17536
rect 37936 17524 37964 17623
rect 38013 17595 38071 17601
rect 38013 17561 38025 17595
rect 38059 17592 38071 17595
rect 38562 17592 38568 17604
rect 38059 17564 38568 17592
rect 38059 17561 38071 17564
rect 38013 17555 38071 17561
rect 38562 17552 38568 17564
rect 38620 17592 38626 17604
rect 38841 17595 38899 17601
rect 38841 17592 38853 17595
rect 38620 17564 38853 17592
rect 38620 17552 38626 17564
rect 38841 17561 38853 17564
rect 38887 17561 38899 17595
rect 43272 17592 43300 17623
rect 43438 17620 43444 17632
rect 43496 17620 43502 17672
rect 43625 17663 43683 17669
rect 43625 17629 43637 17663
rect 43671 17629 43683 17663
rect 43625 17623 43683 17629
rect 43530 17592 43536 17604
rect 43272 17564 43536 17592
rect 38841 17555 38899 17561
rect 43530 17552 43536 17564
rect 43588 17552 43594 17604
rect 43640 17592 43668 17623
rect 43714 17620 43720 17672
rect 43772 17660 43778 17672
rect 43772 17632 43817 17660
rect 43772 17620 43778 17632
rect 44174 17620 44180 17672
rect 44232 17660 44238 17672
rect 44545 17663 44603 17669
rect 44545 17660 44557 17663
rect 44232 17632 44557 17660
rect 44232 17620 44238 17632
rect 44545 17629 44557 17632
rect 44591 17660 44603 17663
rect 45278 17660 45284 17672
rect 44591 17632 45284 17660
rect 44591 17629 44603 17632
rect 44545 17623 44603 17629
rect 45278 17620 45284 17632
rect 45336 17660 45342 17672
rect 45373 17663 45431 17669
rect 45373 17660 45385 17663
rect 45336 17632 45385 17660
rect 45336 17620 45342 17632
rect 45373 17629 45385 17632
rect 45419 17629 45431 17663
rect 45373 17623 45431 17629
rect 45462 17620 45468 17672
rect 45520 17660 45526 17672
rect 45649 17663 45707 17669
rect 45520 17632 45565 17660
rect 45520 17620 45526 17632
rect 45649 17629 45661 17663
rect 45695 17629 45707 17663
rect 45649 17623 45707 17629
rect 45094 17592 45100 17604
rect 43640 17564 45100 17592
rect 45094 17552 45100 17564
rect 45152 17592 45158 17604
rect 45664 17592 45692 17623
rect 45738 17620 45744 17672
rect 45796 17660 45802 17672
rect 46382 17660 46388 17672
rect 45796 17632 45841 17660
rect 46343 17632 46388 17660
rect 45796 17620 45802 17632
rect 46382 17620 46388 17632
rect 46440 17620 46446 17672
rect 46477 17663 46535 17669
rect 46477 17650 46489 17663
rect 46523 17650 46535 17663
rect 46584 17660 46612 17700
rect 46845 17663 46903 17669
rect 46845 17660 46857 17663
rect 46014 17592 46020 17604
rect 45152 17564 46020 17592
rect 45152 17552 45158 17564
rect 46014 17552 46020 17564
rect 46072 17552 46078 17604
rect 46474 17598 46480 17650
rect 46532 17598 46538 17650
rect 46584 17632 46857 17660
rect 46845 17629 46857 17632
rect 46891 17629 46903 17663
rect 47302 17660 47308 17672
rect 46845 17623 46903 17629
rect 46952 17632 47308 17660
rect 46661 17595 46719 17601
rect 46661 17561 46673 17595
rect 46707 17561 46719 17595
rect 46661 17555 46719 17561
rect 46751 17595 46809 17601
rect 46751 17561 46763 17595
rect 46797 17592 46809 17595
rect 46952 17592 46980 17632
rect 47302 17620 47308 17632
rect 47360 17620 47366 17672
rect 47762 17620 47768 17672
rect 47820 17660 47826 17672
rect 49510 17660 49516 17672
rect 47820 17632 49372 17660
rect 49471 17632 49516 17660
rect 47820 17620 47826 17632
rect 47394 17592 47400 17604
rect 46797 17564 46980 17592
rect 47044 17564 47400 17592
rect 46797 17561 46809 17564
rect 46751 17555 46809 17561
rect 36688 17496 37964 17524
rect 36688 17484 36694 17496
rect 38930 17484 38936 17536
rect 38988 17524 38994 17536
rect 39041 17527 39099 17533
rect 39041 17524 39053 17527
rect 38988 17496 39053 17524
rect 38988 17484 38994 17496
rect 39041 17493 39053 17496
rect 39087 17493 39099 17527
rect 39041 17487 39099 17493
rect 39850 17484 39856 17536
rect 39908 17524 39914 17536
rect 40589 17527 40647 17533
rect 40589 17524 40601 17527
rect 39908 17496 40601 17524
rect 39908 17484 39914 17496
rect 40589 17493 40601 17496
rect 40635 17524 40647 17527
rect 40678 17524 40684 17536
rect 40635 17496 40684 17524
rect 40635 17493 40647 17496
rect 40589 17487 40647 17493
rect 40678 17484 40684 17496
rect 40736 17484 40742 17536
rect 42702 17524 42708 17536
rect 42663 17496 42708 17524
rect 42702 17484 42708 17496
rect 42760 17484 42766 17536
rect 46676 17524 46704 17555
rect 46842 17524 46848 17536
rect 46676 17496 46848 17524
rect 46842 17484 46848 17496
rect 46900 17484 46906 17536
rect 47044 17533 47072 17564
rect 47394 17552 47400 17564
rect 47452 17552 47458 17604
rect 48225 17595 48283 17601
rect 48225 17561 48237 17595
rect 48271 17592 48283 17595
rect 48314 17592 48320 17604
rect 48271 17564 48320 17592
rect 48271 17561 48283 17564
rect 48225 17555 48283 17561
rect 48314 17552 48320 17564
rect 48372 17552 48378 17604
rect 49344 17592 49372 17632
rect 49510 17620 49516 17632
rect 49568 17620 49574 17672
rect 49620 17660 49648 17700
rect 49786 17688 49792 17700
rect 49844 17728 49850 17740
rect 50724 17728 50752 17768
rect 52012 17768 52101 17796
rect 52012 17728 52040 17768
rect 52089 17765 52101 17768
rect 52135 17796 52147 17799
rect 52822 17796 52828 17808
rect 52135 17768 52828 17796
rect 52135 17765 52147 17768
rect 52089 17759 52147 17765
rect 52822 17756 52828 17768
rect 52880 17756 52886 17808
rect 53377 17799 53435 17805
rect 53377 17796 53389 17799
rect 53300 17768 53389 17796
rect 52178 17728 52184 17740
rect 49844 17700 50660 17728
rect 50724 17700 52040 17728
rect 52139 17700 52184 17728
rect 49844 17688 49850 17700
rect 50341 17663 50399 17669
rect 50341 17660 50353 17663
rect 49620 17632 50353 17660
rect 50341 17629 50353 17632
rect 50387 17629 50399 17663
rect 50522 17660 50528 17672
rect 50483 17632 50528 17660
rect 50341 17623 50399 17629
rect 50522 17620 50528 17632
rect 50580 17620 50586 17672
rect 50632 17669 50660 17700
rect 52178 17688 52184 17700
rect 52236 17688 52242 17740
rect 52273 17731 52331 17737
rect 52273 17697 52285 17731
rect 52319 17728 52331 17731
rect 52730 17728 52736 17740
rect 52319 17700 52736 17728
rect 52319 17697 52331 17700
rect 52273 17691 52331 17697
rect 52730 17688 52736 17700
rect 52788 17688 52794 17740
rect 50617 17663 50675 17669
rect 50617 17629 50629 17663
rect 50663 17629 50675 17663
rect 50617 17623 50675 17629
rect 50706 17620 50712 17672
rect 50764 17660 50770 17672
rect 50764 17632 50809 17660
rect 50764 17620 50770 17632
rect 51810 17620 51816 17672
rect 51868 17660 51874 17672
rect 51994 17660 52000 17672
rect 51868 17632 52000 17660
rect 51868 17620 51874 17632
rect 51994 17620 52000 17632
rect 52052 17660 52058 17672
rect 52362 17660 52368 17672
rect 52052 17632 52368 17660
rect 52052 17620 52058 17632
rect 52362 17620 52368 17632
rect 52420 17620 52426 17672
rect 52457 17663 52515 17669
rect 52457 17629 52469 17663
rect 52503 17660 52515 17663
rect 53190 17660 53196 17672
rect 52503 17632 53196 17660
rect 52503 17629 52515 17632
rect 52457 17623 52515 17629
rect 53190 17620 53196 17632
rect 53248 17620 53254 17672
rect 53300 17660 53328 17768
rect 53377 17765 53389 17768
rect 53423 17765 53435 17799
rect 53377 17759 53435 17765
rect 55674 17688 55680 17740
rect 55732 17728 55738 17740
rect 55950 17728 55956 17740
rect 55732 17700 55956 17728
rect 55732 17688 55738 17700
rect 55950 17688 55956 17700
rect 56008 17688 56014 17740
rect 56137 17731 56195 17737
rect 56137 17697 56149 17731
rect 56183 17728 56195 17731
rect 56594 17728 56600 17740
rect 56183 17700 56600 17728
rect 56183 17697 56195 17700
rect 56137 17691 56195 17697
rect 56594 17688 56600 17700
rect 56652 17688 56658 17740
rect 53834 17660 53840 17672
rect 53300 17632 53840 17660
rect 53834 17620 53840 17632
rect 53892 17620 53898 17672
rect 54021 17663 54079 17669
rect 54021 17629 54033 17663
rect 54067 17660 54079 17663
rect 54110 17660 54116 17672
rect 54067 17632 54116 17660
rect 54067 17629 54079 17632
rect 54021 17623 54079 17629
rect 54110 17620 54116 17632
rect 54168 17620 54174 17672
rect 55858 17660 55864 17672
rect 55819 17632 55864 17660
rect 55858 17620 55864 17632
rect 55916 17620 55922 17672
rect 50154 17592 50160 17604
rect 49344 17564 50160 17592
rect 50154 17552 50160 17564
rect 50212 17552 50218 17604
rect 50890 17552 50896 17604
rect 50948 17592 50954 17604
rect 53009 17595 53067 17601
rect 53009 17592 53021 17595
rect 50948 17564 53021 17592
rect 50948 17552 50954 17564
rect 53009 17561 53021 17564
rect 53055 17592 53067 17595
rect 53055 17564 54984 17592
rect 53055 17561 53067 17564
rect 53009 17555 53067 17561
rect 54956 17536 54984 17564
rect 47029 17527 47087 17533
rect 47029 17493 47041 17527
rect 47075 17493 47087 17527
rect 47029 17487 47087 17493
rect 47578 17484 47584 17536
rect 47636 17524 47642 17536
rect 48425 17527 48483 17533
rect 48425 17524 48437 17527
rect 47636 17496 48437 17524
rect 47636 17484 47642 17496
rect 48425 17493 48437 17496
rect 48471 17493 48483 17527
rect 48425 17487 48483 17493
rect 48866 17484 48872 17536
rect 48924 17524 48930 17536
rect 49789 17527 49847 17533
rect 49789 17524 49801 17527
rect 48924 17496 49801 17524
rect 48924 17484 48930 17496
rect 49789 17493 49801 17496
rect 49835 17524 49847 17527
rect 51350 17524 51356 17536
rect 49835 17496 51356 17524
rect 49835 17493 49847 17496
rect 49789 17487 49847 17493
rect 51350 17484 51356 17496
rect 51408 17484 51414 17536
rect 51902 17484 51908 17536
rect 51960 17524 51966 17536
rect 53209 17527 53267 17533
rect 53209 17524 53221 17527
rect 51960 17496 53221 17524
rect 51960 17484 51966 17496
rect 53209 17493 53221 17496
rect 53255 17524 53267 17527
rect 54202 17524 54208 17536
rect 53255 17496 54208 17524
rect 53255 17493 53267 17496
rect 53209 17487 53267 17493
rect 54202 17484 54208 17496
rect 54260 17484 54266 17536
rect 54478 17484 54484 17536
rect 54536 17524 54542 17536
rect 54665 17527 54723 17533
rect 54665 17524 54677 17527
rect 54536 17496 54677 17524
rect 54536 17484 54542 17496
rect 54665 17493 54677 17496
rect 54711 17493 54723 17527
rect 54665 17487 54723 17493
rect 54938 17484 54944 17536
rect 54996 17524 55002 17536
rect 56689 17527 56747 17533
rect 56689 17524 56701 17527
rect 54996 17496 56701 17524
rect 54996 17484 55002 17496
rect 56689 17493 56701 17496
rect 56735 17493 56747 17527
rect 56689 17487 56747 17493
rect 57238 17484 57244 17536
rect 57296 17524 57302 17536
rect 57333 17527 57391 17533
rect 57333 17524 57345 17527
rect 57296 17496 57345 17524
rect 57296 17484 57302 17496
rect 57333 17493 57345 17496
rect 57379 17524 57391 17527
rect 57882 17524 57888 17536
rect 57379 17496 57888 17524
rect 57379 17493 57391 17496
rect 57333 17487 57391 17493
rect 57882 17484 57888 17496
rect 57940 17484 57946 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 22465 17323 22523 17329
rect 22465 17320 22477 17323
rect 22152 17292 22477 17320
rect 22152 17280 22158 17292
rect 22465 17289 22477 17292
rect 22511 17289 22523 17323
rect 22465 17283 22523 17289
rect 24762 17280 24768 17332
rect 24820 17320 24826 17332
rect 24949 17323 25007 17329
rect 24949 17320 24961 17323
rect 24820 17292 24961 17320
rect 24820 17280 24826 17292
rect 24949 17289 24961 17292
rect 24995 17289 25007 17323
rect 24949 17283 25007 17289
rect 25498 17280 25504 17332
rect 25556 17320 25562 17332
rect 25593 17323 25651 17329
rect 25593 17320 25605 17323
rect 25556 17292 25605 17320
rect 25556 17280 25562 17292
rect 25593 17289 25605 17292
rect 25639 17289 25651 17323
rect 25593 17283 25651 17289
rect 27706 17280 27712 17332
rect 27764 17320 27770 17332
rect 31202 17320 31208 17332
rect 27764 17292 30972 17320
rect 31163 17292 31208 17320
rect 27764 17280 27770 17292
rect 27801 17255 27859 17261
rect 27801 17221 27813 17255
rect 27847 17252 27859 17255
rect 30282 17252 30288 17264
rect 27847 17224 30288 17252
rect 27847 17221 27859 17224
rect 27801 17215 27859 17221
rect 22554 17184 22560 17196
rect 22515 17156 22560 17184
rect 22554 17144 22560 17156
rect 22612 17144 22618 17196
rect 24026 17144 24032 17196
rect 24084 17184 24090 17196
rect 24581 17187 24639 17193
rect 24581 17184 24593 17187
rect 24084 17156 24593 17184
rect 24084 17144 24090 17156
rect 24581 17153 24593 17156
rect 24627 17184 24639 17187
rect 24854 17184 24860 17196
rect 24627 17156 24860 17184
rect 24627 17153 24639 17156
rect 24581 17147 24639 17153
rect 24854 17144 24860 17156
rect 24912 17144 24918 17196
rect 25409 17187 25467 17193
rect 25409 17153 25421 17187
rect 25455 17153 25467 17187
rect 25409 17147 25467 17153
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17184 26387 17187
rect 26418 17184 26424 17196
rect 26375 17156 26424 17184
rect 26375 17153 26387 17156
rect 26329 17147 26387 17153
rect 23750 17076 23756 17128
rect 23808 17116 23814 17128
rect 24673 17119 24731 17125
rect 24673 17116 24685 17119
rect 23808 17088 24685 17116
rect 23808 17076 23814 17088
rect 24673 17085 24685 17088
rect 24719 17116 24731 17119
rect 25424 17116 25452 17147
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 26513 17187 26571 17193
rect 26513 17153 26525 17187
rect 26559 17184 26571 17187
rect 27816 17184 27844 17215
rect 30282 17212 30288 17224
rect 30340 17212 30346 17264
rect 26559 17156 27844 17184
rect 27985 17187 28043 17193
rect 26559 17153 26571 17156
rect 26513 17147 26571 17153
rect 27985 17153 27997 17187
rect 28031 17184 28043 17187
rect 28074 17184 28080 17196
rect 28031 17156 28080 17184
rect 28031 17153 28043 17156
rect 27985 17147 28043 17153
rect 28074 17144 28080 17156
rect 28132 17144 28138 17196
rect 29086 17144 29092 17196
rect 29144 17184 29150 17196
rect 29181 17187 29239 17193
rect 29181 17184 29193 17187
rect 29144 17156 29193 17184
rect 29144 17144 29150 17156
rect 29181 17153 29193 17156
rect 29227 17153 29239 17187
rect 29181 17147 29239 17153
rect 29273 17187 29331 17193
rect 29273 17153 29285 17187
rect 29319 17153 29331 17187
rect 29273 17147 29331 17153
rect 29457 17187 29515 17193
rect 29457 17153 29469 17187
rect 29503 17184 29515 17187
rect 29917 17187 29975 17193
rect 29917 17184 29929 17187
rect 29503 17156 29929 17184
rect 29503 17153 29515 17156
rect 29457 17147 29515 17153
rect 29917 17153 29929 17156
rect 29963 17153 29975 17187
rect 30558 17184 30564 17196
rect 30519 17156 30564 17184
rect 29917 17147 29975 17153
rect 29288 17116 29316 17147
rect 24719 17088 25452 17116
rect 28644 17088 29316 17116
rect 24719 17085 24731 17088
rect 24673 17079 24731 17085
rect 23566 16940 23572 16992
rect 23624 16980 23630 16992
rect 23845 16983 23903 16989
rect 23845 16980 23857 16983
rect 23624 16952 23857 16980
rect 23624 16940 23630 16952
rect 23845 16949 23857 16952
rect 23891 16949 23903 16983
rect 23845 16943 23903 16949
rect 24765 16983 24823 16989
rect 24765 16949 24777 16983
rect 24811 16980 24823 16983
rect 25682 16980 25688 16992
rect 24811 16952 25688 16980
rect 24811 16949 24823 16952
rect 24765 16943 24823 16949
rect 25682 16940 25688 16952
rect 25740 16940 25746 16992
rect 26234 16940 26240 16992
rect 26292 16980 26298 16992
rect 26513 16983 26571 16989
rect 26513 16980 26525 16983
rect 26292 16952 26525 16980
rect 26292 16940 26298 16952
rect 26513 16949 26525 16952
rect 26559 16949 26571 16983
rect 27614 16980 27620 16992
rect 27575 16952 27620 16980
rect 26513 16943 26571 16949
rect 27614 16940 27620 16952
rect 27672 16940 27678 16992
rect 28442 16940 28448 16992
rect 28500 16980 28506 16992
rect 28644 16989 28672 17088
rect 28994 17008 29000 17060
rect 29052 17048 29058 17060
rect 29472 17048 29500 17147
rect 29932 17116 29960 17147
rect 30558 17144 30564 17156
rect 30616 17144 30622 17196
rect 30650 17144 30656 17196
rect 30708 17184 30714 17196
rect 30944 17193 30972 17292
rect 31202 17280 31208 17292
rect 31260 17280 31266 17332
rect 32677 17323 32735 17329
rect 32677 17289 32689 17323
rect 32723 17320 32735 17323
rect 33134 17320 33140 17332
rect 32723 17292 33140 17320
rect 32723 17289 32735 17292
rect 32677 17283 32735 17289
rect 33134 17280 33140 17292
rect 33192 17280 33198 17332
rect 34054 17320 34060 17332
rect 34015 17292 34060 17320
rect 34054 17280 34060 17292
rect 34112 17280 34118 17332
rect 35253 17323 35311 17329
rect 35253 17289 35265 17323
rect 35299 17320 35311 17323
rect 35526 17320 35532 17332
rect 35299 17292 35532 17320
rect 35299 17289 35311 17292
rect 35253 17283 35311 17289
rect 35526 17280 35532 17292
rect 35584 17280 35590 17332
rect 35618 17280 35624 17332
rect 35676 17320 35682 17332
rect 35713 17323 35771 17329
rect 35713 17320 35725 17323
rect 35676 17292 35725 17320
rect 35676 17280 35682 17292
rect 35713 17289 35725 17292
rect 35759 17289 35771 17323
rect 35713 17283 35771 17289
rect 37274 17280 37280 17332
rect 37332 17320 37338 17332
rect 37461 17323 37519 17329
rect 37461 17320 37473 17323
rect 37332 17292 37473 17320
rect 37332 17280 37338 17292
rect 37461 17289 37473 17292
rect 37507 17289 37519 17323
rect 37461 17283 37519 17289
rect 38562 17280 38568 17332
rect 38620 17320 38626 17332
rect 38841 17323 38899 17329
rect 38841 17320 38853 17323
rect 38620 17292 38853 17320
rect 38620 17280 38626 17292
rect 38841 17289 38853 17292
rect 38887 17289 38899 17323
rect 38841 17283 38899 17289
rect 40221 17323 40279 17329
rect 40221 17289 40233 17323
rect 40267 17320 40279 17323
rect 40865 17323 40923 17329
rect 40865 17320 40877 17323
rect 40267 17292 40877 17320
rect 40267 17289 40279 17292
rect 40221 17283 40279 17289
rect 40865 17289 40877 17292
rect 40911 17320 40923 17323
rect 41138 17320 41144 17332
rect 40911 17292 41144 17320
rect 40911 17289 40923 17292
rect 40865 17283 40923 17289
rect 41138 17280 41144 17292
rect 41196 17280 41202 17332
rect 42981 17323 43039 17329
rect 42981 17289 42993 17323
rect 43027 17320 43039 17323
rect 43438 17320 43444 17332
rect 43027 17292 43444 17320
rect 43027 17289 43039 17292
rect 42981 17283 43039 17289
rect 43438 17280 43444 17292
rect 43496 17280 43502 17332
rect 43530 17280 43536 17332
rect 43588 17320 43594 17332
rect 43809 17323 43867 17329
rect 43809 17320 43821 17323
rect 43588 17292 43821 17320
rect 43588 17280 43594 17292
rect 43809 17289 43821 17292
rect 43855 17289 43867 17323
rect 46106 17320 46112 17332
rect 46067 17292 46112 17320
rect 43809 17283 43867 17289
rect 46106 17280 46112 17292
rect 46164 17280 46170 17332
rect 46382 17280 46388 17332
rect 46440 17320 46446 17332
rect 46753 17323 46811 17329
rect 46753 17320 46765 17323
rect 46440 17292 46765 17320
rect 46440 17280 46446 17292
rect 46753 17289 46765 17292
rect 46799 17289 46811 17323
rect 46753 17283 46811 17289
rect 46842 17280 46848 17332
rect 46900 17320 46906 17332
rect 47118 17320 47124 17332
rect 46900 17292 47124 17320
rect 46900 17280 46906 17292
rect 47118 17280 47124 17292
rect 47176 17280 47182 17332
rect 50341 17323 50399 17329
rect 50341 17289 50353 17323
rect 50387 17320 50399 17323
rect 51442 17320 51448 17332
rect 50387 17292 51448 17320
rect 50387 17289 50399 17292
rect 50341 17283 50399 17289
rect 51442 17280 51448 17292
rect 51500 17280 51506 17332
rect 51537 17323 51595 17329
rect 51537 17289 51549 17323
rect 51583 17320 51595 17323
rect 53006 17320 53012 17332
rect 51583 17292 53012 17320
rect 51583 17289 51595 17292
rect 51537 17283 51595 17289
rect 53006 17280 53012 17292
rect 53064 17280 53070 17332
rect 53926 17320 53932 17332
rect 53887 17292 53932 17320
rect 53926 17280 53932 17292
rect 53984 17280 53990 17332
rect 54481 17323 54539 17329
rect 54481 17289 54493 17323
rect 54527 17320 54539 17323
rect 54570 17320 54576 17332
rect 54527 17292 54576 17320
rect 54527 17289 54539 17292
rect 54481 17283 54539 17289
rect 54570 17280 54576 17292
rect 54628 17280 54634 17332
rect 56410 17320 56416 17332
rect 56371 17292 56416 17320
rect 56410 17280 56416 17292
rect 56468 17280 56474 17332
rect 57422 17320 57428 17332
rect 57383 17292 57428 17320
rect 57422 17280 57428 17292
rect 57480 17280 57486 17332
rect 34793 17255 34851 17261
rect 34793 17252 34805 17255
rect 33796 17224 34805 17252
rect 33796 17196 33824 17224
rect 34793 17221 34805 17224
rect 34839 17252 34851 17255
rect 36081 17255 36139 17261
rect 36081 17252 36093 17255
rect 34839 17224 36093 17252
rect 34839 17221 34851 17224
rect 34793 17215 34851 17221
rect 36081 17221 36093 17224
rect 36127 17221 36139 17255
rect 40678 17252 40684 17264
rect 40639 17224 40684 17252
rect 36081 17215 36139 17221
rect 40678 17212 40684 17224
rect 40736 17212 40742 17264
rect 45646 17212 45652 17264
rect 45704 17252 45710 17264
rect 47765 17255 47823 17261
rect 47765 17252 47777 17255
rect 45704 17224 47777 17252
rect 45704 17212 45710 17224
rect 30745 17187 30803 17193
rect 30745 17184 30757 17187
rect 30708 17156 30757 17184
rect 30708 17144 30714 17156
rect 30745 17153 30757 17156
rect 30791 17153 30803 17187
rect 30745 17147 30803 17153
rect 30837 17187 30895 17193
rect 30837 17153 30849 17187
rect 30883 17153 30895 17187
rect 30837 17147 30895 17153
rect 30929 17187 30987 17193
rect 30929 17153 30941 17187
rect 30975 17153 30987 17187
rect 30929 17147 30987 17153
rect 30466 17116 30472 17128
rect 29932 17088 30472 17116
rect 30466 17076 30472 17088
rect 30524 17076 30530 17128
rect 30852 17116 30880 17147
rect 31018 17144 31024 17196
rect 31076 17184 31082 17196
rect 32493 17187 32551 17193
rect 32493 17184 32505 17187
rect 31076 17156 32505 17184
rect 31076 17144 31082 17156
rect 32493 17153 32505 17156
rect 32539 17153 32551 17187
rect 32493 17147 32551 17153
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17184 33747 17187
rect 33778 17184 33784 17196
rect 33735 17156 33784 17184
rect 33735 17153 33747 17156
rect 33689 17147 33747 17153
rect 33778 17144 33784 17156
rect 33836 17144 33842 17196
rect 33873 17187 33931 17193
rect 33873 17153 33885 17187
rect 33919 17184 33931 17187
rect 34146 17184 34152 17196
rect 33919 17156 34152 17184
rect 33919 17153 33931 17156
rect 33873 17147 33931 17153
rect 31570 17116 31576 17128
rect 30852 17088 31576 17116
rect 31570 17076 31576 17088
rect 31628 17076 31634 17128
rect 32306 17116 32312 17128
rect 32267 17088 32312 17116
rect 32306 17076 32312 17088
rect 32364 17076 32370 17128
rect 32950 17076 32956 17128
rect 33008 17116 33014 17128
rect 33888 17116 33916 17147
rect 34146 17144 34152 17156
rect 34204 17144 34210 17196
rect 34698 17144 34704 17196
rect 34756 17184 34762 17196
rect 34885 17187 34943 17193
rect 34885 17184 34897 17187
rect 34756 17156 34897 17184
rect 34756 17144 34762 17156
rect 34885 17153 34897 17156
rect 34931 17184 34943 17187
rect 36173 17187 36231 17193
rect 36173 17184 36185 17187
rect 34931 17156 36185 17184
rect 34931 17153 34943 17156
rect 34885 17147 34943 17153
rect 36173 17153 36185 17156
rect 36219 17153 36231 17187
rect 37734 17184 37740 17196
rect 37695 17156 37740 17184
rect 36173 17147 36231 17153
rect 37734 17144 37740 17156
rect 37792 17144 37798 17196
rect 38746 17184 38752 17196
rect 38707 17156 38752 17184
rect 38746 17144 38752 17156
rect 38804 17144 38810 17196
rect 38930 17144 38936 17196
rect 38988 17184 38994 17196
rect 39025 17187 39083 17193
rect 39025 17184 39037 17187
rect 38988 17156 39037 17184
rect 38988 17144 38994 17156
rect 39025 17153 39037 17156
rect 39071 17153 39083 17187
rect 39942 17184 39948 17196
rect 39903 17156 39948 17184
rect 39025 17147 39083 17153
rect 39942 17144 39948 17156
rect 40000 17144 40006 17196
rect 40034 17144 40040 17196
rect 40092 17184 40098 17196
rect 40129 17187 40187 17193
rect 40129 17184 40141 17187
rect 40092 17156 40141 17184
rect 40092 17144 40098 17156
rect 40129 17153 40141 17156
rect 40175 17153 40187 17187
rect 40129 17147 40187 17153
rect 40218 17144 40224 17196
rect 40276 17184 40282 17196
rect 42702 17184 42708 17196
rect 40276 17156 40321 17184
rect 42663 17156 42708 17184
rect 40276 17144 40282 17156
rect 42702 17144 42708 17156
rect 42760 17144 42766 17196
rect 43438 17184 43444 17196
rect 43399 17156 43444 17184
rect 43438 17144 43444 17156
rect 43496 17144 43502 17196
rect 43625 17187 43683 17193
rect 43625 17153 43637 17187
rect 43671 17184 43683 17187
rect 43806 17184 43812 17196
rect 43671 17156 43812 17184
rect 43671 17153 43683 17156
rect 43625 17147 43683 17153
rect 34606 17116 34612 17128
rect 33008 17088 33916 17116
rect 34567 17088 34612 17116
rect 33008 17076 33014 17088
rect 34606 17076 34612 17088
rect 34664 17076 34670 17128
rect 36262 17076 36268 17128
rect 36320 17116 36326 17128
rect 37458 17116 37464 17128
rect 36320 17088 36365 17116
rect 37419 17088 37464 17116
rect 36320 17076 36326 17088
rect 37458 17076 37464 17088
rect 37516 17076 37522 17128
rect 42981 17119 43039 17125
rect 42981 17085 42993 17119
rect 43027 17116 43039 17119
rect 43456 17116 43484 17144
rect 43027 17088 43484 17116
rect 43027 17085 43039 17088
rect 42981 17079 43039 17085
rect 29052 17020 29500 17048
rect 29052 17008 29058 17020
rect 30558 17008 30564 17060
rect 30616 17048 30622 17060
rect 32968 17048 32996 17076
rect 30616 17020 32996 17048
rect 30616 17008 30622 17020
rect 36906 17008 36912 17060
rect 36964 17048 36970 17060
rect 38378 17048 38384 17060
rect 36964 17020 38384 17048
rect 36964 17008 36970 17020
rect 38378 17008 38384 17020
rect 38436 17008 38442 17060
rect 39022 17048 39028 17060
rect 38983 17020 39028 17048
rect 39022 17008 39028 17020
rect 39080 17008 39086 17060
rect 42061 17051 42119 17057
rect 42061 17017 42073 17051
rect 42107 17048 42119 17051
rect 43640 17048 43668 17147
rect 43806 17144 43812 17156
rect 43864 17144 43870 17196
rect 44634 17184 44640 17196
rect 44595 17156 44640 17184
rect 44634 17144 44640 17156
rect 44692 17144 44698 17196
rect 44821 17187 44879 17193
rect 44821 17153 44833 17187
rect 44867 17153 44879 17187
rect 45922 17184 45928 17196
rect 45835 17156 45928 17184
rect 44821 17147 44879 17153
rect 44266 17076 44272 17128
rect 44324 17116 44330 17128
rect 44836 17116 44864 17147
rect 45922 17144 45928 17156
rect 45980 17144 45986 17196
rect 46124 17193 46152 17224
rect 47765 17221 47777 17224
rect 47811 17252 47823 17255
rect 48314 17252 48320 17264
rect 47811 17224 48320 17252
rect 47811 17221 47823 17224
rect 47765 17215 47823 17221
rect 48314 17212 48320 17224
rect 48372 17252 48378 17264
rect 49326 17252 49332 17264
rect 48372 17224 49332 17252
rect 48372 17212 48378 17224
rect 49326 17212 49332 17224
rect 49384 17252 49390 17264
rect 49384 17224 49740 17252
rect 49384 17212 49390 17224
rect 46109 17187 46167 17193
rect 46109 17153 46121 17187
rect 46155 17153 46167 17187
rect 46109 17147 46167 17153
rect 46937 17187 46995 17193
rect 46937 17153 46949 17187
rect 46983 17184 46995 17187
rect 47121 17187 47179 17193
rect 46983 17156 47072 17184
rect 46983 17153 46995 17156
rect 46937 17147 46995 17153
rect 44324 17088 44864 17116
rect 45940 17116 45968 17144
rect 45940 17088 46152 17116
rect 44324 17076 44330 17088
rect 46124 17060 46152 17088
rect 42107 17020 43668 17048
rect 44729 17051 44787 17057
rect 42107 17017 42119 17020
rect 42061 17011 42119 17017
rect 44729 17017 44741 17051
rect 44775 17048 44787 17051
rect 45554 17048 45560 17060
rect 44775 17020 45560 17048
rect 44775 17017 44787 17020
rect 44729 17011 44787 17017
rect 45554 17008 45560 17020
rect 45612 17008 45618 17060
rect 46106 17008 46112 17060
rect 46164 17008 46170 17060
rect 47044 17048 47072 17156
rect 47121 17153 47133 17187
rect 47167 17184 47179 17187
rect 48866 17184 48872 17196
rect 47167 17156 48872 17184
rect 47167 17153 47179 17156
rect 47121 17147 47179 17153
rect 48866 17144 48872 17156
rect 48924 17144 48930 17196
rect 48958 17144 48964 17196
rect 49016 17184 49022 17196
rect 49513 17187 49571 17193
rect 49513 17184 49525 17187
rect 49016 17156 49061 17184
rect 49160 17156 49525 17184
rect 49016 17144 49022 17156
rect 47210 17116 47216 17128
rect 47171 17088 47216 17116
rect 47210 17076 47216 17088
rect 47268 17076 47274 17128
rect 48056 17116 48314 17127
rect 48498 17116 48504 17128
rect 47320 17099 48504 17116
rect 47320 17088 48084 17099
rect 48286 17088 48504 17099
rect 47320 17048 47348 17088
rect 48498 17076 48504 17088
rect 48556 17076 48562 17128
rect 49050 17076 49056 17128
rect 49108 17116 49114 17128
rect 49160 17116 49188 17156
rect 49513 17153 49525 17156
rect 49559 17153 49571 17187
rect 49513 17147 49571 17153
rect 49712 17125 49740 17224
rect 50706 17212 50712 17264
rect 50764 17252 50770 17264
rect 52730 17252 52736 17264
rect 50764 17224 52736 17252
rect 50764 17212 50770 17224
rect 50430 17184 50436 17196
rect 50391 17156 50436 17184
rect 50430 17144 50436 17156
rect 50488 17144 50494 17196
rect 51000 17193 51028 17224
rect 52730 17212 52736 17224
rect 52788 17212 52794 17264
rect 52822 17212 52828 17264
rect 52880 17252 52886 17264
rect 52880 17224 53972 17252
rect 52880 17212 52886 17224
rect 53944 17196 53972 17224
rect 54110 17212 54116 17264
rect 54168 17252 54174 17264
rect 54665 17255 54723 17261
rect 54665 17252 54677 17255
rect 54168 17224 54677 17252
rect 54168 17212 54174 17224
rect 54665 17221 54677 17224
rect 54711 17221 54723 17255
rect 54665 17215 54723 17221
rect 50985 17187 51043 17193
rect 50985 17153 50997 17187
rect 51031 17153 51043 17187
rect 50985 17147 51043 17153
rect 51169 17187 51227 17193
rect 51169 17153 51181 17187
rect 51215 17153 51227 17187
rect 51261 17187 51319 17193
rect 51261 17158 51273 17187
rect 51307 17158 51319 17187
rect 51169 17147 51227 17153
rect 49108 17088 49188 17116
rect 49237 17119 49295 17125
rect 49108 17076 49114 17088
rect 49237 17085 49249 17119
rect 49283 17085 49295 17119
rect 49237 17079 49295 17085
rect 49697 17119 49755 17125
rect 49697 17085 49709 17119
rect 49743 17116 49755 17119
rect 50062 17116 50068 17128
rect 49743 17088 50068 17116
rect 49743 17085 49755 17088
rect 49697 17079 49755 17085
rect 47044 17020 47348 17048
rect 48314 17008 48320 17060
rect 48372 17048 48378 17060
rect 49252 17048 49280 17079
rect 50062 17076 50068 17088
rect 50120 17076 50126 17128
rect 51184 17048 51212 17147
rect 51258 17106 51264 17158
rect 51316 17106 51322 17158
rect 51350 17144 51356 17196
rect 51408 17184 51414 17196
rect 51994 17184 52000 17196
rect 51408 17156 51453 17184
rect 51955 17156 52000 17184
rect 51408 17144 51414 17156
rect 51994 17144 52000 17156
rect 52052 17144 52058 17196
rect 53006 17144 53012 17196
rect 53064 17184 53070 17196
rect 53285 17187 53343 17193
rect 53285 17184 53297 17187
rect 53064 17156 53297 17184
rect 53064 17144 53070 17156
rect 53285 17153 53297 17156
rect 53331 17153 53343 17187
rect 53834 17184 53840 17196
rect 53795 17156 53840 17184
rect 53285 17147 53343 17153
rect 53834 17144 53840 17156
rect 53892 17144 53898 17196
rect 53926 17144 53932 17196
rect 53984 17144 53990 17196
rect 54021 17187 54079 17193
rect 54021 17153 54033 17187
rect 54067 17153 54079 17187
rect 54846 17184 54852 17196
rect 54807 17156 54852 17184
rect 54021 17147 54079 17153
rect 51902 17076 51908 17128
rect 51960 17116 51966 17128
rect 52089 17119 52147 17125
rect 52089 17116 52101 17119
rect 51960 17088 52101 17116
rect 51960 17076 51966 17088
rect 52089 17085 52101 17088
rect 52135 17085 52147 17119
rect 52089 17079 52147 17085
rect 52273 17119 52331 17125
rect 52273 17085 52285 17119
rect 52319 17116 52331 17119
rect 52362 17116 52368 17128
rect 52319 17088 52368 17116
rect 52319 17085 52331 17088
rect 52273 17079 52331 17085
rect 52362 17076 52368 17088
rect 52420 17076 52426 17128
rect 53650 17116 53656 17128
rect 53024 17088 53656 17116
rect 52181 17051 52239 17057
rect 52181 17048 52193 17051
rect 48372 17020 49280 17048
rect 50080 17020 51120 17048
rect 51184 17020 52193 17048
rect 48372 17008 48378 17020
rect 28629 16983 28687 16989
rect 28629 16980 28641 16983
rect 28500 16952 28641 16980
rect 28500 16940 28506 16952
rect 28629 16949 28641 16952
rect 28675 16949 28687 16983
rect 29454 16980 29460 16992
rect 29415 16952 29460 16980
rect 28629 16943 28687 16949
rect 29454 16940 29460 16952
rect 29512 16940 29518 16992
rect 37182 16940 37188 16992
rect 37240 16980 37246 16992
rect 37645 16983 37703 16989
rect 37645 16980 37657 16983
rect 37240 16952 37657 16980
rect 37240 16940 37246 16952
rect 37645 16949 37657 16952
rect 37691 16949 37703 16983
rect 40862 16980 40868 16992
rect 40823 16952 40868 16980
rect 37645 16943 37703 16949
rect 40862 16940 40868 16952
rect 40920 16940 40926 16992
rect 41049 16983 41107 16989
rect 41049 16949 41061 16983
rect 41095 16980 41107 16983
rect 41506 16980 41512 16992
rect 41095 16952 41512 16980
rect 41095 16949 41107 16952
rect 41049 16943 41107 16949
rect 41506 16940 41512 16952
rect 41564 16940 41570 16992
rect 42518 16940 42524 16992
rect 42576 16980 42582 16992
rect 42797 16983 42855 16989
rect 42797 16980 42809 16983
rect 42576 16952 42809 16980
rect 42576 16940 42582 16952
rect 42797 16949 42809 16952
rect 42843 16980 42855 16983
rect 43441 16983 43499 16989
rect 43441 16980 43453 16983
rect 42843 16952 43453 16980
rect 42843 16949 42855 16952
rect 42797 16943 42855 16949
rect 43441 16949 43453 16952
rect 43487 16949 43499 16983
rect 43441 16943 43499 16949
rect 45094 16940 45100 16992
rect 45152 16980 45158 16992
rect 45281 16983 45339 16989
rect 45281 16980 45293 16983
rect 45152 16952 45293 16980
rect 45152 16940 45158 16952
rect 45281 16949 45293 16952
rect 45327 16949 45339 16983
rect 45281 16943 45339 16949
rect 45462 16940 45468 16992
rect 45520 16980 45526 16992
rect 50080 16980 50108 17020
rect 45520 16952 50108 16980
rect 45520 16940 45526 16952
rect 50154 16940 50160 16992
rect 50212 16980 50218 16992
rect 50798 16980 50804 16992
rect 50212 16952 50804 16980
rect 50212 16940 50218 16952
rect 50798 16940 50804 16952
rect 50856 16940 50862 16992
rect 51092 16980 51120 17020
rect 52181 17017 52193 17020
rect 52227 17017 52239 17051
rect 52181 17011 52239 17017
rect 51994 16980 52000 16992
rect 51092 16952 52000 16980
rect 51994 16940 52000 16952
rect 52052 16940 52058 16992
rect 52730 16940 52736 16992
rect 52788 16980 52794 16992
rect 53024 16989 53052 17088
rect 53650 17076 53656 17088
rect 53708 17116 53714 17128
rect 54036 17116 54064 17147
rect 54846 17144 54852 17156
rect 54904 17144 54910 17196
rect 55858 17184 55864 17196
rect 55819 17156 55864 17184
rect 55858 17144 55864 17156
rect 55916 17144 55922 17196
rect 55950 17144 55956 17196
rect 56008 17184 56014 17196
rect 56137 17187 56195 17193
rect 56137 17184 56149 17187
rect 56008 17156 56149 17184
rect 56008 17144 56014 17156
rect 56137 17153 56149 17156
rect 56183 17153 56195 17187
rect 56137 17147 56195 17153
rect 56229 17187 56287 17193
rect 56229 17153 56241 17187
rect 56275 17184 56287 17187
rect 56502 17184 56508 17196
rect 56275 17156 56508 17184
rect 56275 17153 56287 17156
rect 56229 17147 56287 17153
rect 56502 17144 56508 17156
rect 56560 17144 56566 17196
rect 54202 17116 54208 17128
rect 53708 17088 54208 17116
rect 53708 17076 53714 17088
rect 54202 17076 54208 17088
rect 54260 17116 54266 17128
rect 54478 17116 54484 17128
rect 54260 17088 54484 17116
rect 54260 17076 54266 17088
rect 54478 17076 54484 17088
rect 54536 17116 54542 17128
rect 56873 17119 56931 17125
rect 56873 17116 56885 17119
rect 54536 17088 56885 17116
rect 54536 17076 54542 17088
rect 56873 17085 56885 17088
rect 56919 17116 56931 17119
rect 57514 17116 57520 17128
rect 56919 17088 57520 17116
rect 56919 17085 56931 17088
rect 56873 17079 56931 17085
rect 57514 17076 57520 17088
rect 57572 17116 57578 17128
rect 58069 17119 58127 17125
rect 58069 17116 58081 17119
rect 57572 17088 58081 17116
rect 57572 17076 57578 17088
rect 58069 17085 58081 17088
rect 58115 17085 58127 17119
rect 58069 17079 58127 17085
rect 55401 17051 55459 17057
rect 55401 17017 55413 17051
rect 55447 17048 55459 17051
rect 55674 17048 55680 17060
rect 55447 17020 55680 17048
rect 55447 17017 55459 17020
rect 55401 17011 55459 17017
rect 55674 17008 55680 17020
rect 55732 17008 55738 17060
rect 53009 16983 53067 16989
rect 53009 16980 53021 16983
rect 52788 16952 53021 16980
rect 52788 16940 52794 16952
rect 53009 16949 53021 16952
rect 53055 16949 53067 16983
rect 53009 16943 53067 16949
rect 55490 16940 55496 16992
rect 55548 16980 55554 16992
rect 55953 16983 56011 16989
rect 55953 16980 55965 16983
rect 55548 16952 55965 16980
rect 55548 16940 55554 16952
rect 55953 16949 55965 16952
rect 55999 16949 56011 16983
rect 55953 16943 56011 16949
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 23750 16736 23756 16788
rect 23808 16776 23814 16788
rect 24029 16779 24087 16785
rect 24029 16776 24041 16779
rect 23808 16748 24041 16776
rect 23808 16736 23814 16748
rect 24029 16745 24041 16748
rect 24075 16745 24087 16779
rect 28994 16776 29000 16788
rect 28955 16748 29000 16776
rect 24029 16739 24087 16745
rect 28994 16736 29000 16748
rect 29052 16736 29058 16788
rect 30926 16736 30932 16788
rect 30984 16776 30990 16788
rect 31205 16779 31263 16785
rect 31205 16776 31217 16779
rect 30984 16748 31217 16776
rect 30984 16736 30990 16748
rect 31205 16745 31217 16748
rect 31251 16745 31263 16779
rect 31205 16739 31263 16745
rect 31570 16736 31576 16788
rect 31628 16776 31634 16788
rect 31628 16748 37136 16776
rect 31628 16736 31634 16748
rect 26510 16708 26516 16720
rect 26471 16680 26516 16708
rect 26510 16668 26516 16680
rect 26568 16668 26574 16720
rect 27893 16711 27951 16717
rect 27893 16677 27905 16711
rect 27939 16708 27951 16711
rect 27982 16708 27988 16720
rect 27939 16680 27988 16708
rect 27939 16677 27951 16680
rect 27893 16671 27951 16677
rect 27982 16668 27988 16680
rect 28040 16668 28046 16720
rect 29181 16711 29239 16717
rect 29181 16677 29193 16711
rect 29227 16708 29239 16711
rect 29730 16708 29736 16720
rect 29227 16680 29736 16708
rect 29227 16677 29239 16680
rect 29181 16671 29239 16677
rect 29730 16668 29736 16680
rect 29788 16708 29794 16720
rect 29788 16680 29960 16708
rect 29788 16668 29794 16680
rect 22094 16600 22100 16652
rect 22152 16640 22158 16652
rect 22281 16643 22339 16649
rect 22281 16640 22293 16643
rect 22152 16612 22293 16640
rect 22152 16600 22158 16612
rect 22281 16609 22293 16612
rect 22327 16609 22339 16643
rect 22281 16603 22339 16609
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16640 22615 16643
rect 23750 16640 23756 16652
rect 22603 16612 23756 16640
rect 22603 16609 22615 16612
rect 22557 16603 22615 16609
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 26234 16640 26240 16652
rect 26195 16612 26240 16640
rect 26234 16600 26240 16612
rect 26292 16600 26298 16652
rect 27614 16640 27620 16652
rect 27575 16612 27620 16640
rect 27614 16600 27620 16612
rect 27672 16600 27678 16652
rect 29932 16649 29960 16680
rect 30282 16668 30288 16720
rect 30340 16708 30346 16720
rect 32306 16708 32312 16720
rect 30340 16680 32312 16708
rect 30340 16668 30346 16680
rect 32306 16668 32312 16680
rect 32364 16668 32370 16720
rect 36725 16711 36783 16717
rect 36725 16677 36737 16711
rect 36771 16708 36783 16711
rect 36906 16708 36912 16720
rect 36771 16680 36912 16708
rect 36771 16677 36783 16680
rect 36725 16671 36783 16677
rect 36906 16668 36912 16680
rect 36964 16668 36970 16720
rect 37108 16717 37136 16748
rect 39316 16748 39804 16776
rect 37093 16711 37151 16717
rect 37093 16677 37105 16711
rect 37139 16677 37151 16711
rect 37093 16671 37151 16677
rect 29917 16643 29975 16649
rect 29917 16609 29929 16643
rect 29963 16609 29975 16643
rect 29917 16603 29975 16609
rect 33134 16600 33140 16652
rect 33192 16640 33198 16652
rect 33321 16643 33379 16649
rect 33321 16640 33333 16643
rect 33192 16612 33333 16640
rect 33192 16600 33198 16612
rect 33321 16609 33333 16612
rect 33367 16609 33379 16643
rect 33321 16603 33379 16609
rect 37001 16643 37059 16649
rect 37001 16609 37013 16643
rect 37047 16609 37059 16643
rect 38378 16640 38384 16652
rect 38339 16612 38384 16640
rect 37001 16603 37059 16609
rect 26142 16572 26148 16584
rect 26103 16544 26148 16572
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26602 16532 26608 16584
rect 26660 16572 26666 16584
rect 27525 16575 27583 16581
rect 27525 16572 27537 16575
rect 26660 16544 27537 16572
rect 26660 16532 26666 16544
rect 27525 16541 27537 16544
rect 27571 16541 27583 16575
rect 27525 16535 27583 16541
rect 29043 16541 29101 16547
rect 29043 16538 29055 16541
rect 23842 16504 23848 16516
rect 23755 16476 23848 16504
rect 23842 16464 23848 16476
rect 23900 16504 23906 16516
rect 24673 16507 24731 16513
rect 24673 16504 24685 16507
rect 23900 16476 24685 16504
rect 23900 16464 23906 16476
rect 24673 16473 24685 16476
rect 24719 16504 24731 16507
rect 24762 16504 24768 16516
rect 24719 16476 24768 16504
rect 24719 16473 24731 16476
rect 24673 16467 24731 16473
rect 24762 16464 24768 16476
rect 24820 16504 24826 16516
rect 25498 16504 25504 16516
rect 24820 16476 25504 16504
rect 24820 16464 24826 16476
rect 25498 16464 25504 16476
rect 25556 16504 25562 16516
rect 28442 16504 28448 16516
rect 25556 16476 28448 16504
rect 25556 16464 25562 16476
rect 28442 16464 28448 16476
rect 28500 16504 28506 16516
rect 28813 16507 28871 16513
rect 28813 16504 28825 16507
rect 28500 16476 28825 16504
rect 28500 16464 28506 16476
rect 28813 16473 28825 16476
rect 28859 16473 28871 16507
rect 29028 16507 29055 16538
rect 29089 16516 29101 16541
rect 29454 16532 29460 16584
rect 29512 16572 29518 16584
rect 30009 16575 30067 16581
rect 30009 16572 30021 16575
rect 29512 16544 30021 16572
rect 29512 16532 29518 16544
rect 30009 16541 30021 16544
rect 30055 16541 30067 16575
rect 30009 16535 30067 16541
rect 30190 16532 30196 16584
rect 30248 16572 30254 16584
rect 30285 16575 30343 16581
rect 30285 16572 30297 16575
rect 30248 16544 30297 16572
rect 30248 16532 30254 16544
rect 30285 16541 30297 16544
rect 30331 16541 30343 16575
rect 30285 16535 30343 16541
rect 30466 16532 30472 16584
rect 30524 16572 30530 16584
rect 31113 16575 31171 16581
rect 31113 16572 31125 16575
rect 30524 16544 31125 16572
rect 30524 16532 30530 16544
rect 31113 16541 31125 16544
rect 31159 16541 31171 16575
rect 31113 16535 31171 16541
rect 31202 16532 31208 16584
rect 31260 16572 31266 16584
rect 31297 16575 31355 16581
rect 31297 16572 31309 16575
rect 31260 16544 31309 16572
rect 31260 16532 31266 16544
rect 31297 16541 31309 16544
rect 31343 16541 31355 16575
rect 31297 16535 31355 16541
rect 31941 16575 31999 16581
rect 31941 16541 31953 16575
rect 31987 16541 31999 16575
rect 31941 16535 31999 16541
rect 29089 16507 29092 16516
rect 29028 16476 29092 16507
rect 28813 16467 28871 16473
rect 29086 16464 29092 16476
rect 29144 16464 29150 16516
rect 31956 16504 31984 16535
rect 33042 16532 33048 16584
rect 33100 16572 33106 16584
rect 33778 16572 33784 16584
rect 33100 16544 33784 16572
rect 33100 16532 33106 16544
rect 33778 16532 33784 16544
rect 33836 16572 33842 16584
rect 33965 16575 34023 16581
rect 33965 16572 33977 16575
rect 33836 16544 33977 16572
rect 33836 16532 33842 16544
rect 33965 16541 33977 16544
rect 34011 16541 34023 16575
rect 34146 16572 34152 16584
rect 34107 16544 34152 16572
rect 33965 16535 34023 16541
rect 34146 16532 34152 16544
rect 34204 16532 34210 16584
rect 36630 16532 36636 16584
rect 36688 16572 36694 16584
rect 36909 16575 36967 16581
rect 36909 16572 36921 16575
rect 36688 16544 36921 16572
rect 36688 16532 36694 16544
rect 36909 16541 36921 16544
rect 36955 16541 36967 16575
rect 36909 16535 36967 16541
rect 32950 16504 32956 16516
rect 30116 16476 32956 16504
rect 26234 16396 26240 16448
rect 26292 16436 26298 16448
rect 26510 16436 26516 16448
rect 26292 16408 26516 16436
rect 26292 16396 26298 16408
rect 26510 16396 26516 16408
rect 26568 16436 26574 16448
rect 27154 16436 27160 16448
rect 26568 16408 27160 16436
rect 26568 16396 26574 16408
rect 27154 16396 27160 16408
rect 27212 16436 27218 16448
rect 30116 16436 30144 16476
rect 32950 16464 32956 16476
rect 33008 16504 33014 16516
rect 33229 16507 33287 16513
rect 33229 16504 33241 16507
rect 33008 16476 33241 16504
rect 33008 16464 33014 16476
rect 33229 16473 33241 16476
rect 33275 16504 33287 16507
rect 34698 16504 34704 16516
rect 33275 16476 34704 16504
rect 33275 16473 33287 16476
rect 33229 16467 33287 16473
rect 34698 16464 34704 16476
rect 34756 16464 34762 16516
rect 30282 16436 30288 16448
rect 27212 16408 30144 16436
rect 30243 16408 30288 16436
rect 27212 16396 27218 16408
rect 30282 16396 30288 16408
rect 30340 16396 30346 16448
rect 31294 16396 31300 16448
rect 31352 16436 31358 16448
rect 31849 16439 31907 16445
rect 31849 16436 31861 16439
rect 31352 16408 31861 16436
rect 31352 16396 31358 16408
rect 31849 16405 31861 16408
rect 31895 16405 31907 16439
rect 32766 16436 32772 16448
rect 32727 16408 32772 16436
rect 31849 16399 31907 16405
rect 32766 16396 32772 16408
rect 32824 16396 32830 16448
rect 33042 16396 33048 16448
rect 33100 16436 33106 16448
rect 33137 16439 33195 16445
rect 33137 16436 33149 16439
rect 33100 16408 33149 16436
rect 33100 16396 33106 16408
rect 33137 16405 33149 16408
rect 33183 16405 33195 16439
rect 33137 16399 33195 16405
rect 34149 16439 34207 16445
rect 34149 16405 34161 16439
rect 34195 16436 34207 16439
rect 34514 16436 34520 16448
rect 34195 16408 34520 16436
rect 34195 16405 34207 16408
rect 34149 16399 34207 16405
rect 34514 16396 34520 16408
rect 34572 16396 34578 16448
rect 37016 16436 37044 16603
rect 38378 16600 38384 16612
rect 38436 16600 38442 16652
rect 39316 16649 39344 16748
rect 39408 16680 39712 16708
rect 39301 16643 39359 16649
rect 39301 16640 39313 16643
rect 38580 16612 39313 16640
rect 38580 16584 38608 16612
rect 39301 16609 39313 16612
rect 39347 16609 39359 16643
rect 39301 16603 39359 16609
rect 37185 16575 37243 16581
rect 37185 16541 37197 16575
rect 37231 16541 37243 16575
rect 37366 16572 37372 16584
rect 37327 16544 37372 16572
rect 37185 16535 37243 16541
rect 37200 16504 37228 16535
rect 37366 16532 37372 16544
rect 37424 16532 37430 16584
rect 38010 16532 38016 16584
rect 38068 16572 38074 16584
rect 38289 16575 38347 16581
rect 38289 16572 38301 16575
rect 38068 16544 38301 16572
rect 38068 16532 38074 16544
rect 38289 16541 38301 16544
rect 38335 16572 38347 16575
rect 38562 16572 38568 16584
rect 38335 16544 38568 16572
rect 38335 16541 38347 16544
rect 38289 16535 38347 16541
rect 38562 16532 38568 16544
rect 38620 16532 38626 16584
rect 38746 16532 38752 16584
rect 38804 16572 38810 16584
rect 39117 16575 39175 16581
rect 39117 16572 39129 16575
rect 38804 16544 39129 16572
rect 38804 16532 38810 16544
rect 39117 16541 39129 16544
rect 39163 16572 39175 16575
rect 39408 16572 39436 16680
rect 39163 16544 39436 16572
rect 39163 16541 39175 16544
rect 39117 16535 39175 16541
rect 39482 16532 39488 16584
rect 39540 16572 39546 16584
rect 39684 16572 39712 16680
rect 39776 16640 39804 16748
rect 40218 16736 40224 16788
rect 40276 16776 40282 16788
rect 40497 16779 40555 16785
rect 40497 16776 40509 16779
rect 40276 16748 40509 16776
rect 40276 16736 40282 16748
rect 40497 16745 40509 16748
rect 40543 16745 40555 16779
rect 40497 16739 40555 16745
rect 42702 16736 42708 16788
rect 42760 16776 42766 16788
rect 44085 16779 44143 16785
rect 44085 16776 44097 16779
rect 42760 16748 44097 16776
rect 42760 16736 42766 16748
rect 44085 16745 44097 16748
rect 44131 16776 44143 16779
rect 45462 16776 45468 16788
rect 44131 16748 45468 16776
rect 44131 16745 44143 16748
rect 44085 16739 44143 16745
rect 45462 16736 45468 16748
rect 45520 16736 45526 16788
rect 47854 16736 47860 16788
rect 47912 16776 47918 16788
rect 52270 16776 52276 16788
rect 47912 16748 48452 16776
rect 47912 16736 47918 16748
rect 48424 16720 48452 16748
rect 51184 16748 52276 16776
rect 47504 16680 47808 16708
rect 39776 16612 40172 16640
rect 40144 16581 40172 16612
rect 40037 16575 40095 16581
rect 40037 16572 40049 16575
rect 39540 16544 39585 16572
rect 39684 16544 40049 16572
rect 39540 16532 39546 16544
rect 40037 16541 40049 16544
rect 40083 16541 40095 16575
rect 40037 16535 40095 16541
rect 40129 16575 40187 16581
rect 40129 16541 40141 16575
rect 40175 16541 40187 16575
rect 40310 16572 40316 16584
rect 40271 16544 40316 16572
rect 40129 16535 40187 16541
rect 40310 16532 40316 16544
rect 40368 16532 40374 16584
rect 41506 16572 41512 16584
rect 41467 16544 41512 16572
rect 41506 16532 41512 16544
rect 41564 16532 41570 16584
rect 41966 16572 41972 16584
rect 41927 16544 41972 16572
rect 41966 16532 41972 16544
rect 42024 16532 42030 16584
rect 44726 16532 44732 16584
rect 44784 16572 44790 16584
rect 45833 16575 45891 16581
rect 45833 16572 45845 16575
rect 44784 16544 45845 16572
rect 44784 16532 44790 16544
rect 45833 16541 45845 16544
rect 45879 16541 45891 16575
rect 46106 16572 46112 16584
rect 46067 16544 46112 16572
rect 45833 16535 45891 16541
rect 46106 16532 46112 16544
rect 46164 16532 46170 16584
rect 46201 16575 46259 16581
rect 46201 16541 46213 16575
rect 46247 16541 46259 16575
rect 46474 16572 46480 16584
rect 46435 16544 46480 16572
rect 46201 16535 46259 16541
rect 37458 16504 37464 16516
rect 37200 16476 37464 16504
rect 37458 16464 37464 16476
rect 37516 16504 37522 16516
rect 39209 16507 39267 16513
rect 37516 16476 38148 16504
rect 37516 16464 37522 16476
rect 38120 16448 38148 16476
rect 39209 16473 39221 16507
rect 39255 16504 39267 16507
rect 40328 16504 40356 16532
rect 39255 16476 40356 16504
rect 39255 16473 39267 16476
rect 39209 16467 39267 16473
rect 42058 16464 42064 16516
rect 42116 16504 42122 16516
rect 43806 16504 43812 16516
rect 42116 16476 42366 16504
rect 43767 16476 43812 16504
rect 42116 16464 42122 16476
rect 43806 16464 43812 16476
rect 43864 16464 43870 16516
rect 45370 16504 45376 16516
rect 45331 16476 45376 16504
rect 45370 16464 45376 16476
rect 45428 16464 45434 16516
rect 37274 16436 37280 16448
rect 37016 16408 37280 16436
rect 37274 16396 37280 16408
rect 37332 16396 37338 16448
rect 37826 16436 37832 16448
rect 37787 16408 37832 16436
rect 37826 16396 37832 16408
rect 37884 16396 37890 16448
rect 38102 16396 38108 16448
rect 38160 16436 38166 16448
rect 38197 16439 38255 16445
rect 38197 16436 38209 16439
rect 38160 16408 38209 16436
rect 38160 16396 38166 16408
rect 38197 16405 38209 16408
rect 38243 16405 38255 16439
rect 38197 16399 38255 16405
rect 39393 16439 39451 16445
rect 39393 16405 39405 16439
rect 39439 16436 39451 16439
rect 40034 16436 40040 16448
rect 39439 16408 40040 16436
rect 39439 16405 39451 16408
rect 39393 16399 39451 16405
rect 40034 16396 40040 16408
rect 40092 16396 40098 16448
rect 46216 16436 46244 16535
rect 46474 16532 46480 16544
rect 46532 16532 46538 16584
rect 46661 16575 46719 16581
rect 46661 16541 46673 16575
rect 46707 16572 46719 16575
rect 46842 16572 46848 16584
rect 46707 16544 46848 16572
rect 46707 16541 46719 16544
rect 46661 16535 46719 16541
rect 46842 16532 46848 16544
rect 46900 16572 46906 16584
rect 47394 16572 47400 16584
rect 46900 16544 47400 16572
rect 46900 16532 46906 16544
rect 47394 16532 47400 16544
rect 47452 16532 47458 16584
rect 46750 16464 46756 16516
rect 46808 16504 46814 16516
rect 47504 16504 47532 16680
rect 47780 16640 47808 16680
rect 48038 16668 48044 16720
rect 48096 16668 48102 16720
rect 48406 16668 48412 16720
rect 48464 16708 48470 16720
rect 48961 16711 49019 16717
rect 48961 16708 48973 16711
rect 48464 16680 48973 16708
rect 48464 16668 48470 16680
rect 48961 16677 48973 16680
rect 49007 16677 49019 16711
rect 48961 16671 49019 16677
rect 50798 16668 50804 16720
rect 50856 16708 50862 16720
rect 51184 16708 51212 16748
rect 52270 16736 52276 16748
rect 52328 16776 52334 16788
rect 52457 16779 52515 16785
rect 52457 16776 52469 16779
rect 52328 16748 52469 16776
rect 52328 16736 52334 16748
rect 52457 16745 52469 16748
rect 52503 16745 52515 16779
rect 52457 16739 52515 16745
rect 52825 16779 52883 16785
rect 52825 16745 52837 16779
rect 52871 16776 52883 16779
rect 53466 16776 53472 16788
rect 52871 16748 53472 16776
rect 52871 16745 52883 16748
rect 52825 16739 52883 16745
rect 53466 16736 53472 16748
rect 53524 16736 53530 16788
rect 53742 16776 53748 16788
rect 53703 16748 53748 16776
rect 53742 16736 53748 16748
rect 53800 16736 53806 16788
rect 54481 16779 54539 16785
rect 54481 16745 54493 16779
rect 54527 16776 54539 16779
rect 54846 16776 54852 16788
rect 54527 16748 54852 16776
rect 54527 16745 54539 16748
rect 54481 16739 54539 16745
rect 54846 16736 54852 16748
rect 54904 16736 54910 16788
rect 56042 16776 56048 16788
rect 56003 16748 56048 16776
rect 56042 16736 56048 16748
rect 56100 16736 56106 16788
rect 56594 16776 56600 16788
rect 56555 16748 56600 16776
rect 56594 16736 56600 16748
rect 56652 16736 56658 16788
rect 53006 16708 53012 16720
rect 50856 16680 51212 16708
rect 51460 16680 53012 16708
rect 50856 16668 50862 16680
rect 48056 16640 48084 16668
rect 48133 16643 48191 16649
rect 48133 16640 48145 16643
rect 47780 16612 47992 16640
rect 48056 16612 48145 16640
rect 47765 16575 47823 16581
rect 47765 16541 47777 16575
rect 47811 16572 47823 16575
rect 47854 16572 47860 16584
rect 47811 16544 47860 16572
rect 47811 16541 47823 16544
rect 47765 16535 47823 16541
rect 47854 16532 47860 16544
rect 47912 16532 47918 16584
rect 47964 16581 47992 16612
rect 48133 16609 48145 16612
rect 48179 16609 48191 16643
rect 48133 16603 48191 16609
rect 48774 16600 48780 16652
rect 48832 16640 48838 16652
rect 51460 16640 51488 16680
rect 53006 16668 53012 16680
rect 53064 16668 53070 16720
rect 48832 16612 49188 16640
rect 48832 16600 48838 16612
rect 49160 16581 49188 16612
rect 50540 16612 51488 16640
rect 50540 16584 50568 16612
rect 47949 16575 48007 16581
rect 47949 16541 47961 16575
rect 47995 16541 48007 16575
rect 47949 16535 48007 16541
rect 48225 16575 48283 16581
rect 48225 16541 48237 16575
rect 48271 16541 48283 16575
rect 48225 16535 48283 16541
rect 48501 16575 48559 16581
rect 48501 16541 48513 16575
rect 48547 16572 48559 16575
rect 49145 16575 49203 16581
rect 48547 16544 48820 16572
rect 48547 16541 48559 16544
rect 48501 16535 48559 16541
rect 46808 16476 47532 16504
rect 48240 16504 48268 16535
rect 48792 16516 48820 16544
rect 49145 16541 49157 16575
rect 49191 16572 49203 16575
rect 50062 16572 50068 16584
rect 49191 16544 50068 16572
rect 49191 16541 49203 16544
rect 49145 16535 49203 16541
rect 50062 16532 50068 16544
rect 50120 16532 50126 16584
rect 50522 16572 50528 16584
rect 50483 16544 50528 16572
rect 50522 16532 50528 16544
rect 50580 16532 50586 16584
rect 50709 16575 50767 16581
rect 50709 16541 50721 16575
rect 50755 16572 50767 16575
rect 50798 16572 50804 16584
rect 50755 16544 50804 16572
rect 50755 16541 50767 16544
rect 50709 16535 50767 16541
rect 50798 16532 50804 16544
rect 50856 16532 50862 16584
rect 51350 16572 51356 16584
rect 51311 16544 51356 16572
rect 51350 16532 51356 16544
rect 51408 16532 51414 16584
rect 51460 16581 51488 16612
rect 52365 16643 52423 16649
rect 52365 16609 52377 16643
rect 52411 16640 52423 16643
rect 52546 16640 52552 16652
rect 52411 16612 52552 16640
rect 52411 16609 52423 16612
rect 52365 16603 52423 16609
rect 52546 16600 52552 16612
rect 52604 16600 52610 16652
rect 53098 16600 53104 16652
rect 53156 16640 53162 16652
rect 53156 16612 53604 16640
rect 53156 16600 53162 16612
rect 51445 16575 51503 16581
rect 51445 16541 51457 16575
rect 51491 16541 51503 16575
rect 51445 16535 51503 16541
rect 51721 16575 51779 16581
rect 51721 16541 51733 16575
rect 51767 16541 51779 16575
rect 52638 16572 52644 16584
rect 52599 16544 52644 16572
rect 51721 16535 51779 16541
rect 48240 16476 48531 16504
rect 46808 16464 46814 16476
rect 48503 16448 48531 16476
rect 48774 16464 48780 16516
rect 48832 16464 48838 16516
rect 49329 16507 49387 16513
rect 49329 16473 49341 16507
rect 49375 16504 49387 16507
rect 49602 16504 49608 16516
rect 49375 16476 49608 16504
rect 49375 16473 49387 16476
rect 49329 16467 49387 16473
rect 49602 16464 49608 16476
rect 49660 16464 49666 16516
rect 50617 16507 50675 16513
rect 50617 16473 50629 16507
rect 50663 16504 50675 16507
rect 50663 16476 51396 16504
rect 50663 16473 50675 16476
rect 50617 16467 50675 16473
rect 48268 16436 48274 16448
rect 46216 16408 48274 16436
rect 48268 16396 48274 16408
rect 48326 16396 48332 16448
rect 48498 16396 48504 16448
rect 48556 16396 48562 16448
rect 50982 16396 50988 16448
rect 51040 16436 51046 16448
rect 51169 16439 51227 16445
rect 51169 16436 51181 16439
rect 51040 16408 51181 16436
rect 51040 16396 51046 16408
rect 51169 16405 51181 16408
rect 51215 16405 51227 16439
rect 51368 16436 51396 16476
rect 51534 16464 51540 16516
rect 51592 16504 51598 16516
rect 51592 16476 51637 16504
rect 51592 16464 51598 16476
rect 51736 16436 51764 16535
rect 52638 16532 52644 16544
rect 52696 16532 52702 16584
rect 53285 16575 53343 16581
rect 53285 16541 53297 16575
rect 53331 16572 53343 16575
rect 53374 16572 53380 16584
rect 53331 16544 53380 16572
rect 53331 16541 53343 16544
rect 53285 16535 53343 16541
rect 53374 16532 53380 16544
rect 53432 16532 53438 16584
rect 53576 16581 53604 16612
rect 53834 16600 53840 16652
rect 53892 16640 53898 16652
rect 56502 16640 56508 16652
rect 53892 16612 54800 16640
rect 53892 16600 53898 16612
rect 53561 16575 53619 16581
rect 53561 16541 53573 16575
rect 53607 16572 53619 16575
rect 54662 16572 54668 16584
rect 53607 16544 54524 16572
rect 54623 16544 54668 16572
rect 53607 16541 53619 16544
rect 53561 16535 53619 16541
rect 54496 16516 54524 16544
rect 54662 16532 54668 16544
rect 54720 16532 54726 16584
rect 54772 16581 54800 16612
rect 55784 16612 56088 16640
rect 56463 16612 56508 16640
rect 54757 16575 54815 16581
rect 54757 16541 54769 16575
rect 54803 16572 54815 16575
rect 55030 16572 55036 16584
rect 54803 16544 55036 16572
rect 54803 16541 54815 16544
rect 54757 16535 54815 16541
rect 55030 16532 55036 16544
rect 55088 16532 55094 16584
rect 55490 16572 55496 16584
rect 55451 16544 55496 16572
rect 55490 16532 55496 16544
rect 55548 16532 55554 16584
rect 55582 16532 55588 16584
rect 55640 16572 55646 16584
rect 55784 16581 55812 16612
rect 55769 16575 55827 16581
rect 55640 16544 55685 16572
rect 55640 16532 55646 16544
rect 55769 16541 55781 16575
rect 55815 16541 55827 16575
rect 55769 16535 55827 16541
rect 55861 16575 55919 16581
rect 55861 16541 55873 16575
rect 55907 16541 55919 16575
rect 56060 16572 56088 16612
rect 56502 16600 56508 16612
rect 56560 16600 56566 16652
rect 56689 16643 56747 16649
rect 56689 16609 56701 16643
rect 56735 16609 56747 16643
rect 56689 16603 56747 16609
rect 56704 16572 56732 16603
rect 56060 16544 56732 16572
rect 55861 16535 55919 16541
rect 52270 16464 52276 16516
rect 52328 16504 52334 16516
rect 53190 16504 53196 16516
rect 52328 16476 53196 16504
rect 52328 16464 52334 16476
rect 53190 16464 53196 16476
rect 53248 16464 53254 16516
rect 54478 16504 54484 16516
rect 54439 16476 54484 16504
rect 54478 16464 54484 16476
rect 54536 16464 54542 16516
rect 54680 16504 54708 16532
rect 55784 16504 55812 16535
rect 54680 16476 55812 16504
rect 55876 16504 55904 16535
rect 56778 16532 56784 16584
rect 56836 16572 56842 16584
rect 56836 16544 56881 16572
rect 56836 16532 56842 16544
rect 56686 16504 56692 16516
rect 55876 16476 56692 16504
rect 51368 16408 51764 16436
rect 51169 16399 51227 16405
rect 52546 16396 52552 16448
rect 52604 16436 52610 16448
rect 53377 16439 53435 16445
rect 53377 16436 53389 16439
rect 52604 16408 53389 16436
rect 52604 16396 52610 16408
rect 53377 16405 53389 16408
rect 53423 16405 53435 16439
rect 53377 16399 53435 16405
rect 53742 16396 53748 16448
rect 53800 16436 53806 16448
rect 55876 16436 55904 16476
rect 56686 16464 56692 16476
rect 56744 16504 56750 16516
rect 56962 16504 56968 16516
rect 56744 16476 56968 16504
rect 56744 16464 56750 16476
rect 56962 16464 56968 16476
rect 57020 16464 57026 16516
rect 53800 16408 55904 16436
rect 53800 16396 53806 16408
rect 56594 16396 56600 16448
rect 56652 16436 56658 16448
rect 57241 16439 57299 16445
rect 57241 16436 57253 16439
rect 56652 16408 57253 16436
rect 56652 16396 56658 16408
rect 57241 16405 57253 16408
rect 57287 16405 57299 16439
rect 57882 16436 57888 16448
rect 57843 16408 57888 16436
rect 57241 16399 57299 16405
rect 57882 16396 57888 16408
rect 57940 16396 57946 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 22094 16232 22100 16244
rect 22020 16204 22100 16232
rect 22020 16105 22048 16204
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 23566 16232 23572 16244
rect 22296 16204 23572 16232
rect 22296 16173 22324 16204
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 23750 16232 23756 16244
rect 23711 16204 23756 16232
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 25498 16232 25504 16244
rect 25459 16204 25504 16232
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 26142 16192 26148 16244
rect 26200 16232 26206 16244
rect 26602 16232 26608 16244
rect 26200 16204 26464 16232
rect 26563 16204 26608 16232
rect 26200 16192 26206 16204
rect 22281 16167 22339 16173
rect 22281 16133 22293 16167
rect 22327 16133 22339 16167
rect 23842 16164 23848 16176
rect 23506 16136 23848 16164
rect 22281 16127 22339 16133
rect 23842 16124 23848 16136
rect 23900 16124 23906 16176
rect 26436 16164 26464 16204
rect 26602 16192 26608 16204
rect 26660 16192 26666 16244
rect 28994 16192 29000 16244
rect 29052 16232 29058 16244
rect 29181 16235 29239 16241
rect 29181 16232 29193 16235
rect 29052 16204 29193 16232
rect 29052 16192 29058 16204
rect 29181 16201 29193 16204
rect 29227 16201 29239 16235
rect 29181 16195 29239 16201
rect 30101 16235 30159 16241
rect 30101 16201 30113 16235
rect 30147 16232 30159 16235
rect 30558 16232 30564 16244
rect 30147 16204 30564 16232
rect 30147 16201 30159 16204
rect 30101 16195 30159 16201
rect 30558 16192 30564 16204
rect 30616 16192 30622 16244
rect 31573 16235 31631 16241
rect 31573 16201 31585 16235
rect 31619 16232 31631 16235
rect 33042 16232 33048 16244
rect 31619 16204 33048 16232
rect 31619 16201 31631 16204
rect 31573 16195 31631 16201
rect 33042 16192 33048 16204
rect 33100 16192 33106 16244
rect 33229 16235 33287 16241
rect 33229 16201 33241 16235
rect 33275 16232 33287 16235
rect 33686 16232 33692 16244
rect 33275 16204 33692 16232
rect 33275 16201 33287 16204
rect 33229 16195 33287 16201
rect 33686 16192 33692 16204
rect 33744 16192 33750 16244
rect 34333 16235 34391 16241
rect 34333 16201 34345 16235
rect 34379 16232 34391 16235
rect 34422 16232 34428 16244
rect 34379 16204 34428 16232
rect 34379 16201 34391 16204
rect 34333 16195 34391 16201
rect 34422 16192 34428 16204
rect 34480 16192 34486 16244
rect 34698 16232 34704 16244
rect 34659 16204 34704 16232
rect 34698 16192 34704 16204
rect 34756 16192 34762 16244
rect 36814 16232 36820 16244
rect 36775 16204 36820 16232
rect 36814 16192 36820 16204
rect 36872 16192 36878 16244
rect 38102 16232 38108 16244
rect 38063 16204 38108 16232
rect 38102 16192 38108 16204
rect 38160 16192 38166 16244
rect 40218 16192 40224 16244
rect 40276 16232 40282 16244
rect 40313 16235 40371 16241
rect 40313 16232 40325 16235
rect 40276 16204 40325 16232
rect 40276 16192 40282 16204
rect 40313 16201 40325 16204
rect 40359 16201 40371 16235
rect 40313 16195 40371 16201
rect 40681 16235 40739 16241
rect 40681 16201 40693 16235
rect 40727 16232 40739 16235
rect 40862 16232 40868 16244
rect 40727 16204 40868 16232
rect 40727 16201 40739 16204
rect 40681 16195 40739 16201
rect 40862 16192 40868 16204
rect 40920 16192 40926 16244
rect 41138 16232 41144 16244
rect 41099 16204 41144 16232
rect 41138 16192 41144 16204
rect 41196 16192 41202 16244
rect 41414 16192 41420 16244
rect 41472 16232 41478 16244
rect 41785 16235 41843 16241
rect 41785 16232 41797 16235
rect 41472 16204 41797 16232
rect 41472 16192 41478 16204
rect 41785 16201 41797 16204
rect 41831 16201 41843 16235
rect 42794 16232 42800 16244
rect 42707 16204 42800 16232
rect 41785 16195 41843 16201
rect 42794 16192 42800 16204
rect 42852 16232 42858 16244
rect 43806 16232 43812 16244
rect 42852 16204 43812 16232
rect 42852 16192 42858 16204
rect 43806 16192 43812 16204
rect 43864 16192 43870 16244
rect 44726 16232 44732 16244
rect 44687 16204 44732 16232
rect 44726 16192 44732 16204
rect 44784 16192 44790 16244
rect 46198 16232 46204 16244
rect 46159 16204 46204 16232
rect 46198 16192 46204 16204
rect 46256 16192 46262 16244
rect 46753 16235 46811 16241
rect 46753 16201 46765 16235
rect 46799 16201 46811 16235
rect 46753 16195 46811 16201
rect 27617 16167 27675 16173
rect 27617 16164 27629 16167
rect 26436 16136 27629 16164
rect 27617 16133 27629 16136
rect 27663 16164 27675 16167
rect 30466 16164 30472 16176
rect 27663 16136 30472 16164
rect 27663 16133 27675 16136
rect 27617 16127 27675 16133
rect 30466 16124 30472 16136
rect 30524 16124 30530 16176
rect 31202 16124 31208 16176
rect 31260 16164 31266 16176
rect 33060 16164 33088 16192
rect 34793 16167 34851 16173
rect 34793 16164 34805 16167
rect 31260 16136 31754 16164
rect 33060 16136 34805 16164
rect 31260 16124 31266 16136
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 26050 16096 26056 16108
rect 24627 16068 26056 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 26050 16056 26056 16068
rect 26108 16056 26114 16108
rect 26418 16096 26424 16108
rect 26379 16068 26424 16096
rect 26418 16056 26424 16068
rect 26476 16056 26482 16108
rect 27430 16096 27436 16108
rect 27391 16068 27436 16096
rect 27430 16056 27436 16068
rect 27488 16056 27494 16108
rect 29730 16096 29736 16108
rect 29691 16068 29736 16096
rect 29730 16056 29736 16068
rect 29788 16056 29794 16108
rect 29914 16096 29920 16108
rect 29875 16068 29920 16096
rect 29914 16056 29920 16068
rect 29972 16096 29978 16108
rect 30190 16096 30196 16108
rect 29972 16068 30196 16096
rect 29972 16056 29978 16068
rect 30190 16056 30196 16068
rect 30248 16056 30254 16108
rect 31018 16096 31024 16108
rect 30979 16068 31024 16096
rect 31018 16056 31024 16068
rect 31076 16056 31082 16108
rect 31113 16099 31171 16105
rect 31113 16065 31125 16099
rect 31159 16065 31171 16099
rect 31294 16096 31300 16108
rect 31255 16068 31300 16096
rect 31113 16059 31171 16065
rect 24673 16031 24731 16037
rect 24673 15997 24685 16031
rect 24719 15997 24731 16031
rect 24673 15991 24731 15997
rect 24949 16031 25007 16037
rect 24949 15997 24961 16031
rect 24995 16028 25007 16031
rect 25038 16028 25044 16040
rect 24995 16000 25044 16028
rect 24995 15997 25007 16000
rect 24949 15991 25007 15997
rect 24688 15960 24716 15991
rect 25038 15988 25044 16000
rect 25096 15988 25102 16040
rect 26142 16028 26148 16040
rect 26103 16000 26148 16028
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 26237 16031 26295 16037
rect 26237 15997 26249 16031
rect 26283 15997 26295 16031
rect 26237 15991 26295 15997
rect 26252 15960 26280 15991
rect 26326 15988 26332 16040
rect 26384 16028 26390 16040
rect 27154 16028 27160 16040
rect 26384 16000 26429 16028
rect 27115 16000 27160 16028
rect 26384 15988 26390 16000
rect 27154 15988 27160 16000
rect 27212 15988 27218 16040
rect 31128 16028 31156 16059
rect 31294 16056 31300 16068
rect 31352 16056 31358 16108
rect 31386 16056 31392 16108
rect 31444 16096 31450 16108
rect 31726 16096 31754 16136
rect 34793 16133 34805 16136
rect 34839 16164 34851 16167
rect 42981 16167 43039 16173
rect 34839 16136 35756 16164
rect 34839 16133 34851 16136
rect 34793 16127 34851 16133
rect 32861 16099 32919 16105
rect 32861 16096 32873 16099
rect 31444 16068 31489 16096
rect 31726 16068 32873 16096
rect 31444 16056 31450 16068
rect 32861 16065 32873 16068
rect 32907 16065 32919 16099
rect 32861 16059 32919 16065
rect 32953 16099 33011 16105
rect 32953 16065 32965 16099
rect 32999 16096 33011 16099
rect 33410 16096 33416 16108
rect 32999 16068 33416 16096
rect 32999 16065 33011 16068
rect 32953 16059 33011 16065
rect 33410 16056 33416 16068
rect 33468 16056 33474 16108
rect 35728 16105 35756 16136
rect 35820 16136 36952 16164
rect 35713 16099 35771 16105
rect 35713 16065 35725 16099
rect 35759 16065 35771 16099
rect 35713 16059 35771 16065
rect 32766 16028 32772 16040
rect 31128 16000 32772 16028
rect 32766 15988 32772 16000
rect 32824 15988 32830 16040
rect 33045 16031 33103 16037
rect 33045 15997 33057 16031
rect 33091 16028 33103 16031
rect 33318 16028 33324 16040
rect 33091 16000 33324 16028
rect 33091 15997 33103 16000
rect 33045 15991 33103 15997
rect 33318 15988 33324 16000
rect 33376 15988 33382 16040
rect 34977 16031 35035 16037
rect 34977 15997 34989 16031
rect 35023 16028 35035 16031
rect 35434 16028 35440 16040
rect 35023 16000 35440 16028
rect 35023 15997 35035 16000
rect 34977 15991 35035 15997
rect 35434 15988 35440 16000
rect 35492 15988 35498 16040
rect 35618 16028 35624 16040
rect 35579 16000 35624 16028
rect 35618 15988 35624 16000
rect 35676 15988 35682 16040
rect 26970 15960 26976 15972
rect 24688 15932 25544 15960
rect 26252 15932 26976 15960
rect 25516 15892 25544 15932
rect 26970 15920 26976 15932
rect 27028 15920 27034 15972
rect 27890 15920 27896 15972
rect 27948 15960 27954 15972
rect 28169 15963 28227 15969
rect 28169 15960 28181 15963
rect 27948 15932 28181 15960
rect 27948 15920 27954 15932
rect 28169 15929 28181 15932
rect 28215 15960 28227 15963
rect 31110 15960 31116 15972
rect 28215 15932 31116 15960
rect 28215 15929 28227 15932
rect 28169 15923 28227 15929
rect 31110 15920 31116 15932
rect 31168 15920 31174 15972
rect 32490 15920 32496 15972
rect 32548 15960 32554 15972
rect 35820 15960 35848 16136
rect 36722 16096 36728 16108
rect 36683 16068 36728 16096
rect 36722 16056 36728 16068
rect 36780 16056 36786 16108
rect 36924 16105 36952 16136
rect 42981 16133 42993 16167
rect 43027 16164 43039 16167
rect 44361 16167 44419 16173
rect 44361 16164 44373 16167
rect 43027 16136 44373 16164
rect 43027 16133 43039 16136
rect 42981 16127 43039 16133
rect 36909 16099 36967 16105
rect 36909 16065 36921 16099
rect 36955 16096 36967 16099
rect 37642 16096 37648 16108
rect 36955 16068 37648 16096
rect 36955 16065 36967 16068
rect 36909 16059 36967 16065
rect 37642 16056 37648 16068
rect 37700 16056 37706 16108
rect 38010 16096 38016 16108
rect 37971 16068 38016 16096
rect 38010 16056 38016 16068
rect 38068 16056 38074 16108
rect 38197 16099 38255 16105
rect 38197 16065 38209 16099
rect 38243 16096 38255 16099
rect 38746 16096 38752 16108
rect 38243 16068 38752 16096
rect 38243 16065 38255 16068
rect 38197 16059 38255 16065
rect 38746 16056 38752 16068
rect 38804 16056 38810 16108
rect 40034 16056 40040 16108
rect 40092 16096 40098 16108
rect 40221 16099 40279 16105
rect 40221 16096 40233 16099
rect 40092 16068 40233 16096
rect 40092 16056 40098 16068
rect 40221 16065 40233 16068
rect 40267 16065 40279 16099
rect 40221 16059 40279 16065
rect 40497 16099 40555 16105
rect 40497 16065 40509 16099
rect 40543 16065 40555 16099
rect 41506 16096 41512 16108
rect 41467 16068 41512 16096
rect 40497 16059 40555 16065
rect 39942 16028 39948 16040
rect 36096 16000 39948 16028
rect 36096 15969 36124 16000
rect 39942 15988 39948 16000
rect 40000 16028 40006 16040
rect 40512 16028 40540 16059
rect 41506 16056 41512 16068
rect 41564 16056 41570 16108
rect 41601 16099 41659 16105
rect 41601 16065 41613 16099
rect 41647 16096 41659 16099
rect 41966 16096 41972 16108
rect 41647 16068 41972 16096
rect 41647 16065 41659 16068
rect 41601 16059 41659 16065
rect 41966 16056 41972 16068
rect 42024 16056 42030 16108
rect 42702 16096 42708 16108
rect 42663 16068 42708 16096
rect 42702 16056 42708 16068
rect 42760 16056 42766 16108
rect 43732 16105 43760 16136
rect 44361 16133 44373 16136
rect 44407 16164 44419 16167
rect 45186 16164 45192 16176
rect 44407 16136 45192 16164
rect 44407 16133 44419 16136
rect 44361 16127 44419 16133
rect 45186 16124 45192 16136
rect 45244 16124 45250 16176
rect 46768 16164 46796 16195
rect 47210 16192 47216 16244
rect 47268 16232 47274 16244
rect 48498 16232 48504 16244
rect 47268 16204 47992 16232
rect 48459 16204 48504 16232
rect 47268 16192 47274 16204
rect 47854 16164 47860 16176
rect 45756 16136 47860 16164
rect 45756 16108 45784 16136
rect 47854 16124 47860 16136
rect 47912 16124 47918 16176
rect 47964 16164 47992 16204
rect 48498 16192 48504 16204
rect 48556 16192 48562 16244
rect 49234 16192 49240 16244
rect 49292 16232 49298 16244
rect 49513 16235 49571 16241
rect 49513 16232 49525 16235
rect 49292 16204 49525 16232
rect 49292 16192 49298 16204
rect 49513 16201 49525 16204
rect 49559 16201 49571 16235
rect 49513 16195 49571 16201
rect 49528 16164 49556 16195
rect 49970 16192 49976 16244
rect 50028 16232 50034 16244
rect 50157 16235 50215 16241
rect 50157 16232 50169 16235
rect 50028 16204 50169 16232
rect 50028 16192 50034 16204
rect 50157 16201 50169 16204
rect 50203 16201 50215 16235
rect 50157 16195 50215 16201
rect 50798 16192 50804 16244
rect 50856 16232 50862 16244
rect 50982 16232 50988 16244
rect 50856 16204 50988 16232
rect 50856 16192 50862 16204
rect 50982 16192 50988 16204
rect 51040 16192 51046 16244
rect 51534 16192 51540 16244
rect 51592 16232 51598 16244
rect 51721 16235 51779 16241
rect 51721 16232 51733 16235
rect 51592 16204 51733 16232
rect 51592 16192 51598 16204
rect 51721 16201 51733 16204
rect 51767 16201 51779 16235
rect 51721 16195 51779 16201
rect 53653 16235 53711 16241
rect 53653 16201 53665 16235
rect 53699 16232 53711 16235
rect 54110 16232 54116 16244
rect 53699 16204 54116 16232
rect 53699 16201 53711 16204
rect 53653 16195 53711 16201
rect 54110 16192 54116 16204
rect 54168 16192 54174 16244
rect 54478 16192 54484 16244
rect 54536 16232 54542 16244
rect 55125 16235 55183 16241
rect 55125 16232 55137 16235
rect 54536 16204 55137 16232
rect 54536 16192 54542 16204
rect 55125 16201 55137 16204
rect 55171 16232 55183 16235
rect 55674 16232 55680 16244
rect 55171 16204 55680 16232
rect 55171 16201 55183 16204
rect 55125 16195 55183 16201
rect 55674 16192 55680 16204
rect 55732 16192 55738 16244
rect 56045 16235 56103 16241
rect 56045 16201 56057 16235
rect 56091 16232 56103 16235
rect 56502 16232 56508 16244
rect 56091 16204 56508 16232
rect 56091 16201 56103 16204
rect 56045 16195 56103 16201
rect 56502 16192 56508 16204
rect 56560 16192 56566 16244
rect 47964 16136 48912 16164
rect 49528 16136 51120 16164
rect 43533 16099 43591 16105
rect 43533 16065 43545 16099
rect 43579 16065 43591 16099
rect 43533 16059 43591 16065
rect 43717 16099 43775 16105
rect 43717 16065 43729 16099
rect 43763 16065 43775 16099
rect 43717 16059 43775 16065
rect 44545 16099 44603 16105
rect 44545 16065 44557 16099
rect 44591 16065 44603 16099
rect 45554 16096 45560 16108
rect 45515 16068 45560 16096
rect 44545 16059 44603 16065
rect 40000 16000 40540 16028
rect 40000 15988 40006 16000
rect 42518 15988 42524 16040
rect 42576 16028 42582 16040
rect 43548 16028 43576 16059
rect 42576 16000 43576 16028
rect 42576 15988 42582 16000
rect 44082 15988 44088 16040
rect 44140 16028 44146 16040
rect 44450 16028 44456 16040
rect 44140 16000 44456 16028
rect 44140 15988 44146 16000
rect 44450 15988 44456 16000
rect 44508 16028 44514 16040
rect 44560 16028 44588 16059
rect 45554 16056 45560 16068
rect 45612 16056 45618 16108
rect 45738 16096 45744 16108
rect 45699 16068 45744 16096
rect 45738 16056 45744 16068
rect 45796 16056 45802 16108
rect 45925 16099 45983 16105
rect 45925 16065 45937 16099
rect 45971 16096 45983 16099
rect 46014 16096 46020 16108
rect 45971 16068 46020 16096
rect 45971 16065 45983 16068
rect 45925 16059 45983 16065
rect 46014 16056 46020 16068
rect 46072 16056 46078 16108
rect 46109 16099 46167 16105
rect 46109 16065 46121 16099
rect 46155 16065 46167 16099
rect 46109 16059 46167 16065
rect 45830 16028 45836 16040
rect 44508 16000 44588 16028
rect 45791 16000 45836 16028
rect 44508 15988 44514 16000
rect 45830 15988 45836 16000
rect 45888 15988 45894 16040
rect 46124 16028 46152 16059
rect 46198 16056 46204 16108
rect 46256 16096 46262 16108
rect 46753 16099 46811 16105
rect 46753 16096 46765 16099
rect 46256 16068 46765 16096
rect 46256 16056 46262 16068
rect 46753 16065 46765 16068
rect 46799 16094 46811 16099
rect 46842 16094 46848 16108
rect 46799 16066 46848 16094
rect 46799 16065 46811 16066
rect 46753 16059 46811 16065
rect 46842 16056 46848 16066
rect 46900 16056 46906 16108
rect 46937 16099 46995 16105
rect 46937 16065 46949 16099
rect 46983 16065 46995 16099
rect 46937 16059 46995 16065
rect 46658 16028 46664 16040
rect 46124 16000 46664 16028
rect 46658 15988 46664 16000
rect 46716 15988 46722 16040
rect 46952 16028 46980 16059
rect 47394 16056 47400 16108
rect 47452 16096 47458 16108
rect 47765 16099 47823 16105
rect 47765 16096 47777 16099
rect 47452 16068 47777 16096
rect 47452 16056 47458 16068
rect 47765 16065 47777 16068
rect 47811 16065 47823 16099
rect 47765 16059 47823 16065
rect 47949 16099 48007 16105
rect 47949 16065 47961 16099
rect 47995 16096 48007 16099
rect 48130 16096 48136 16108
rect 47995 16068 48136 16096
rect 47995 16065 48007 16068
rect 47949 16059 48007 16065
rect 48130 16056 48136 16068
rect 48188 16056 48194 16108
rect 48682 16096 48688 16108
rect 48643 16068 48688 16096
rect 48682 16056 48688 16068
rect 48740 16056 48746 16108
rect 48884 16105 48912 16136
rect 48869 16099 48927 16105
rect 48869 16065 48881 16099
rect 48915 16096 48927 16099
rect 50154 16096 50160 16108
rect 48915 16068 50160 16096
rect 48915 16065 48927 16068
rect 48869 16059 48927 16065
rect 50154 16056 50160 16068
rect 50212 16056 50218 16108
rect 50341 16099 50399 16105
rect 50341 16065 50353 16099
rect 50387 16096 50399 16099
rect 50430 16096 50436 16108
rect 50387 16068 50436 16096
rect 50387 16065 50399 16068
rect 50341 16059 50399 16065
rect 46886 16000 46980 16028
rect 32548 15932 35848 15960
rect 36081 15963 36139 15969
rect 32548 15920 32554 15932
rect 36081 15929 36093 15963
rect 36127 15929 36139 15963
rect 43622 15960 43628 15972
rect 43583 15932 43628 15960
rect 36081 15923 36139 15929
rect 43622 15920 43628 15932
rect 43680 15920 43686 15972
rect 46750 15960 46756 15972
rect 45480 15932 46756 15960
rect 26326 15892 26332 15904
rect 25516 15864 26332 15892
rect 26326 15852 26332 15864
rect 26384 15892 26390 15904
rect 27249 15895 27307 15901
rect 27249 15892 27261 15895
rect 26384 15864 27261 15892
rect 26384 15852 26390 15864
rect 27249 15861 27261 15864
rect 27295 15861 27307 15895
rect 27249 15855 27307 15861
rect 28442 15852 28448 15904
rect 28500 15892 28506 15904
rect 28629 15895 28687 15901
rect 28629 15892 28641 15895
rect 28500 15864 28641 15892
rect 28500 15852 28506 15864
rect 28629 15861 28641 15864
rect 28675 15861 28687 15895
rect 28629 15855 28687 15861
rect 29454 15852 29460 15904
rect 29512 15892 29518 15904
rect 29733 15895 29791 15901
rect 29733 15892 29745 15895
rect 29512 15864 29745 15892
rect 29512 15852 29518 15864
rect 29733 15861 29745 15864
rect 29779 15861 29791 15895
rect 29733 15855 29791 15861
rect 37826 15852 37832 15904
rect 37884 15892 37890 15904
rect 38749 15895 38807 15901
rect 38749 15892 38761 15895
rect 37884 15864 38761 15892
rect 37884 15852 37890 15864
rect 38749 15861 38761 15864
rect 38795 15892 38807 15895
rect 41598 15892 41604 15904
rect 38795 15864 41604 15892
rect 38795 15861 38807 15864
rect 38749 15855 38807 15861
rect 41598 15852 41604 15864
rect 41656 15852 41662 15904
rect 42981 15895 43039 15901
rect 42981 15861 42993 15895
rect 43027 15892 43039 15895
rect 45480 15892 45508 15932
rect 46750 15920 46756 15932
rect 46808 15920 46814 15972
rect 43027 15864 45508 15892
rect 43027 15861 43039 15864
rect 42981 15855 43039 15861
rect 46106 15852 46112 15904
rect 46164 15892 46170 15904
rect 46886 15892 46914 16000
rect 47026 15988 47032 16040
rect 47084 16028 47090 16040
rect 48777 16031 48835 16037
rect 48777 16028 48789 16031
rect 47084 16000 48789 16028
rect 47084 15988 47090 16000
rect 48777 15997 48789 16000
rect 48823 15997 48835 16031
rect 48777 15991 48835 15997
rect 47946 15960 47952 15972
rect 47907 15932 47952 15960
rect 47946 15920 47952 15932
rect 48004 15920 48010 15972
rect 48792 15960 48820 15991
rect 48958 15988 48964 16040
rect 49016 16028 49022 16040
rect 49016 16000 49061 16028
rect 49016 15988 49022 16000
rect 49970 15988 49976 16040
rect 50028 16028 50034 16040
rect 50356 16028 50384 16059
rect 50430 16056 50436 16068
rect 50488 16056 50494 16108
rect 50614 16096 50620 16108
rect 50575 16068 50620 16096
rect 50614 16056 50620 16068
rect 50672 16056 50678 16108
rect 50798 16096 50804 16108
rect 50759 16068 50804 16096
rect 50798 16056 50804 16068
rect 50856 16056 50862 16108
rect 51092 16096 51120 16136
rect 51166 16124 51172 16176
rect 51224 16164 51230 16176
rect 51261 16167 51319 16173
rect 51261 16164 51273 16167
rect 51224 16136 51273 16164
rect 51224 16124 51230 16136
rect 51261 16133 51273 16136
rect 51307 16133 51319 16167
rect 51261 16127 51319 16133
rect 51092 16068 51488 16096
rect 51350 16028 51356 16040
rect 50028 16000 50384 16028
rect 51311 16000 51356 16028
rect 50028 15988 50034 16000
rect 51350 15988 51356 16000
rect 51408 15988 51414 16040
rect 51460 16028 51488 16068
rect 51534 16056 51540 16108
rect 51592 16096 51598 16108
rect 51994 16096 52000 16108
rect 51592 16068 52000 16096
rect 51592 16056 51598 16068
rect 51994 16056 52000 16068
rect 52052 16096 52058 16108
rect 52181 16099 52239 16105
rect 52181 16096 52193 16099
rect 52052 16068 52193 16096
rect 52052 16056 52058 16068
rect 52181 16065 52193 16068
rect 52227 16065 52239 16099
rect 53834 16096 53840 16108
rect 53795 16068 53840 16096
rect 52181 16059 52239 16065
rect 53834 16056 53840 16068
rect 53892 16056 53898 16108
rect 54021 16099 54079 16105
rect 54021 16065 54033 16099
rect 54067 16096 54079 16099
rect 54849 16099 54907 16105
rect 54067 16068 54340 16096
rect 54067 16065 54079 16068
rect 54021 16059 54079 16065
rect 53742 16028 53748 16040
rect 51460 16000 53748 16028
rect 53742 15988 53748 16000
rect 53800 15988 53806 16040
rect 53929 16031 53987 16037
rect 53929 15997 53941 16031
rect 53975 15997 53987 16031
rect 53929 15991 53987 15997
rect 54113 16031 54171 16037
rect 54113 15997 54125 16031
rect 54159 16028 54171 16031
rect 54202 16028 54208 16040
rect 54159 16000 54208 16028
rect 54159 15997 54171 16000
rect 54113 15991 54171 15997
rect 49418 15960 49424 15972
rect 48792 15932 49424 15960
rect 49418 15920 49424 15932
rect 49476 15920 49482 15972
rect 49694 15920 49700 15972
rect 49752 15960 49758 15972
rect 50433 15963 50491 15969
rect 50433 15960 50445 15963
rect 49752 15932 50445 15960
rect 49752 15920 49758 15932
rect 50433 15929 50445 15932
rect 50479 15929 50491 15963
rect 50433 15923 50491 15929
rect 50525 15963 50583 15969
rect 50525 15929 50537 15963
rect 50571 15929 50583 15963
rect 50525 15923 50583 15929
rect 48958 15892 48964 15904
rect 46164 15864 48964 15892
rect 46164 15852 46170 15864
rect 48958 15852 48964 15864
rect 49016 15852 49022 15904
rect 50246 15852 50252 15904
rect 50304 15892 50310 15904
rect 50540 15892 50568 15923
rect 51074 15920 51080 15972
rect 51132 15960 51138 15972
rect 53944 15960 53972 15991
rect 54202 15988 54208 16000
rect 54260 15988 54266 16040
rect 54312 16028 54340 16068
rect 54849 16065 54861 16099
rect 54895 16096 54907 16099
rect 55214 16096 55220 16108
rect 54895 16068 55220 16096
rect 54895 16065 54907 16068
rect 54849 16059 54907 16065
rect 55214 16056 55220 16068
rect 55272 16056 55278 16108
rect 55582 16056 55588 16108
rect 55640 16096 55646 16108
rect 55953 16099 56011 16105
rect 55953 16096 55965 16099
rect 55640 16068 55965 16096
rect 55640 16056 55646 16068
rect 55953 16065 55965 16068
rect 55999 16065 56011 16099
rect 55953 16059 56011 16065
rect 56137 16099 56195 16105
rect 56137 16065 56149 16099
rect 56183 16065 56195 16099
rect 56137 16059 56195 16065
rect 54312 16000 54892 16028
rect 54864 15972 54892 16000
rect 55490 15988 55496 16040
rect 55548 16028 55554 16040
rect 56152 16028 56180 16059
rect 55548 16000 56180 16028
rect 55548 15988 55554 16000
rect 54478 15960 54484 15972
rect 51132 15932 51304 15960
rect 53944 15932 54484 15960
rect 51132 15920 51138 15932
rect 51276 15901 51304 15932
rect 54478 15920 54484 15932
rect 54536 15920 54542 15972
rect 54846 15920 54852 15972
rect 54904 15960 54910 15972
rect 58069 15963 58127 15969
rect 58069 15960 58081 15963
rect 54904 15932 58081 15960
rect 54904 15920 54910 15932
rect 58069 15929 58081 15932
rect 58115 15929 58127 15963
rect 58069 15923 58127 15929
rect 50304 15864 50568 15892
rect 51261 15895 51319 15901
rect 50304 15852 50310 15864
rect 51261 15861 51273 15895
rect 51307 15861 51319 15895
rect 51261 15855 51319 15861
rect 51442 15852 51448 15904
rect 51500 15892 51506 15904
rect 53009 15895 53067 15901
rect 53009 15892 53021 15895
rect 51500 15864 53021 15892
rect 51500 15852 51506 15864
rect 53009 15861 53021 15864
rect 53055 15892 53067 15895
rect 55122 15892 55128 15904
rect 53055 15864 55128 15892
rect 53055 15861 53067 15864
rect 53009 15855 53067 15861
rect 55122 15852 55128 15864
rect 55180 15852 55186 15904
rect 56594 15892 56600 15904
rect 56555 15864 56600 15892
rect 56594 15852 56600 15864
rect 56652 15852 56658 15904
rect 57146 15892 57152 15904
rect 57107 15864 57152 15892
rect 57146 15852 57152 15864
rect 57204 15852 57210 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 23566 15648 23572 15700
rect 23624 15688 23630 15700
rect 24946 15688 24952 15700
rect 23624 15660 24952 15688
rect 23624 15648 23630 15660
rect 24946 15648 24952 15660
rect 25004 15688 25010 15700
rect 25406 15688 25412 15700
rect 25004 15660 25412 15688
rect 25004 15648 25010 15660
rect 25406 15648 25412 15660
rect 25464 15648 25470 15700
rect 26050 15648 26056 15700
rect 26108 15688 26114 15700
rect 26605 15691 26663 15697
rect 26605 15688 26617 15691
rect 26108 15660 26617 15688
rect 26108 15648 26114 15660
rect 26605 15657 26617 15660
rect 26651 15688 26663 15691
rect 27430 15688 27436 15700
rect 26651 15660 27436 15688
rect 26651 15657 26663 15660
rect 26605 15651 26663 15657
rect 27430 15648 27436 15660
rect 27488 15648 27494 15700
rect 28074 15648 28080 15700
rect 28132 15688 28138 15700
rect 30834 15688 30840 15700
rect 28132 15660 30840 15688
rect 28132 15648 28138 15660
rect 30834 15648 30840 15660
rect 30892 15648 30898 15700
rect 31021 15691 31079 15697
rect 31021 15657 31033 15691
rect 31067 15688 31079 15691
rect 31202 15688 31208 15700
rect 31067 15660 31208 15688
rect 31067 15657 31079 15660
rect 31021 15651 31079 15657
rect 31202 15648 31208 15660
rect 31260 15648 31266 15700
rect 32766 15648 32772 15700
rect 32824 15688 32830 15700
rect 32953 15691 33011 15697
rect 32953 15688 32965 15691
rect 32824 15660 32965 15688
rect 32824 15648 32830 15660
rect 32953 15657 32965 15660
rect 32999 15657 33011 15691
rect 35618 15688 35624 15700
rect 35579 15660 35624 15688
rect 32953 15651 33011 15657
rect 35618 15648 35624 15660
rect 35676 15648 35682 15700
rect 36081 15691 36139 15697
rect 36081 15657 36093 15691
rect 36127 15688 36139 15691
rect 36262 15688 36268 15700
rect 36127 15660 36268 15688
rect 36127 15657 36139 15660
rect 36081 15651 36139 15657
rect 36262 15648 36268 15660
rect 36320 15648 36326 15700
rect 37642 15688 37648 15700
rect 37603 15660 37648 15688
rect 37642 15648 37648 15660
rect 37700 15648 37706 15700
rect 38470 15688 38476 15700
rect 38431 15660 38476 15688
rect 38470 15648 38476 15660
rect 38528 15648 38534 15700
rect 41969 15691 42027 15697
rect 41969 15657 41981 15691
rect 42015 15688 42027 15691
rect 45738 15688 45744 15700
rect 42015 15660 45744 15688
rect 42015 15657 42027 15660
rect 41969 15651 42027 15657
rect 45738 15648 45744 15660
rect 45796 15648 45802 15700
rect 45830 15648 45836 15700
rect 45888 15688 45894 15700
rect 46109 15691 46167 15697
rect 46109 15688 46121 15691
rect 45888 15660 46121 15688
rect 45888 15648 45894 15660
rect 46109 15657 46121 15660
rect 46155 15657 46167 15691
rect 47394 15688 47400 15700
rect 46109 15651 46167 15657
rect 46308 15660 47400 15688
rect 24026 15580 24032 15632
rect 24084 15620 24090 15632
rect 24765 15623 24823 15629
rect 24765 15620 24777 15623
rect 24084 15592 24777 15620
rect 24084 15580 24090 15592
rect 24765 15589 24777 15592
rect 24811 15620 24823 15623
rect 26510 15620 26516 15632
rect 24811 15592 26516 15620
rect 24811 15589 24823 15592
rect 24765 15583 24823 15589
rect 26510 15580 26516 15592
rect 26568 15580 26574 15632
rect 27890 15620 27896 15632
rect 27851 15592 27896 15620
rect 27890 15580 27896 15592
rect 27948 15580 27954 15632
rect 27985 15623 28043 15629
rect 27985 15589 27997 15623
rect 28031 15620 28043 15623
rect 28810 15620 28816 15632
rect 28031 15592 28816 15620
rect 28031 15589 28043 15592
rect 27985 15583 28043 15589
rect 28810 15580 28816 15592
rect 28868 15580 28874 15632
rect 29914 15620 29920 15632
rect 28920 15592 29920 15620
rect 21821 15555 21879 15561
rect 21821 15521 21833 15555
rect 21867 15552 21879 15555
rect 22554 15552 22560 15564
rect 21867 15524 22094 15552
rect 22467 15524 22560 15552
rect 21867 15521 21879 15524
rect 21821 15515 21879 15521
rect 22066 15416 22094 15524
rect 22480 15493 22508 15524
rect 22554 15512 22560 15524
rect 22612 15552 22618 15564
rect 24302 15552 24308 15564
rect 22612 15524 24308 15552
rect 22612 15512 22618 15524
rect 24302 15512 24308 15524
rect 24360 15552 24366 15564
rect 28920 15552 28948 15592
rect 29914 15580 29920 15592
rect 29972 15580 29978 15632
rect 32493 15623 32551 15629
rect 32493 15589 32505 15623
rect 32539 15620 32551 15623
rect 36722 15620 36728 15632
rect 32539 15592 36728 15620
rect 32539 15589 32551 15592
rect 32493 15583 32551 15589
rect 36722 15580 36728 15592
rect 36780 15580 36786 15632
rect 42521 15623 42579 15629
rect 42521 15589 42533 15623
rect 42567 15620 42579 15623
rect 42794 15620 42800 15632
rect 42567 15592 42800 15620
rect 42567 15589 42579 15592
rect 42521 15583 42579 15589
rect 42794 15580 42800 15592
rect 42852 15580 42858 15632
rect 43349 15623 43407 15629
rect 43349 15589 43361 15623
rect 43395 15620 43407 15623
rect 44174 15620 44180 15632
rect 43395 15592 44180 15620
rect 43395 15589 43407 15592
rect 43349 15583 43407 15589
rect 44174 15580 44180 15592
rect 44232 15580 44238 15632
rect 44269 15623 44327 15629
rect 44269 15589 44281 15623
rect 44315 15620 44327 15623
rect 44358 15620 44364 15632
rect 44315 15592 44364 15620
rect 44315 15589 44327 15592
rect 44269 15583 44327 15589
rect 44358 15580 44364 15592
rect 44416 15580 44422 15632
rect 44818 15580 44824 15632
rect 44876 15620 44882 15632
rect 46308 15620 46336 15660
rect 47394 15648 47400 15660
rect 47452 15648 47458 15700
rect 47964 15660 48314 15688
rect 47964 15632 47992 15660
rect 44876 15592 46336 15620
rect 44876 15580 44882 15592
rect 29822 15552 29828 15564
rect 24360 15524 28948 15552
rect 29783 15524 29828 15552
rect 24360 15512 24366 15524
rect 29822 15512 29828 15524
rect 29880 15512 29886 15564
rect 30285 15555 30343 15561
rect 30285 15521 30297 15555
rect 30331 15552 30343 15555
rect 35161 15555 35219 15561
rect 30331 15524 35112 15552
rect 30331 15521 30343 15524
rect 30285 15515 30343 15521
rect 22465 15487 22523 15493
rect 22465 15453 22477 15487
rect 22511 15453 22523 15487
rect 22465 15447 22523 15453
rect 22649 15487 22707 15493
rect 22649 15453 22661 15487
rect 22695 15484 22707 15487
rect 22830 15484 22836 15496
rect 22695 15456 22836 15484
rect 22695 15453 22707 15456
rect 22649 15447 22707 15453
rect 22664 15416 22692 15447
rect 22830 15444 22836 15456
rect 22888 15444 22894 15496
rect 23566 15484 23572 15496
rect 23527 15456 23572 15484
rect 23566 15444 23572 15456
rect 23624 15444 23630 15496
rect 23750 15444 23756 15496
rect 23808 15484 23814 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 23808 15456 24593 15484
rect 23808 15444 23814 15456
rect 24581 15453 24593 15456
rect 24627 15484 24639 15487
rect 26053 15487 26111 15493
rect 26053 15484 26065 15487
rect 24627 15456 26065 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 26053 15453 26065 15456
rect 26099 15453 26111 15487
rect 26053 15447 26111 15453
rect 26145 15487 26203 15493
rect 26145 15453 26157 15487
rect 26191 15453 26203 15487
rect 26145 15447 26203 15453
rect 22066 15388 22692 15416
rect 26160 15416 26188 15447
rect 26234 15444 26240 15496
rect 26292 15484 26298 15496
rect 26329 15487 26387 15493
rect 26329 15484 26341 15487
rect 26292 15456 26341 15484
rect 26292 15444 26298 15456
rect 26329 15453 26341 15456
rect 26375 15453 26387 15487
rect 26329 15447 26387 15453
rect 26421 15487 26479 15493
rect 26421 15453 26433 15487
rect 26467 15484 26479 15487
rect 27982 15484 27988 15496
rect 26467 15456 27988 15484
rect 26467 15453 26479 15456
rect 26421 15447 26479 15453
rect 27982 15444 27988 15456
rect 28040 15444 28046 15496
rect 28534 15444 28540 15496
rect 28592 15444 28598 15496
rect 28718 15484 28724 15496
rect 28679 15456 28724 15484
rect 28718 15444 28724 15456
rect 28776 15444 28782 15496
rect 28813 15487 28871 15493
rect 28813 15453 28825 15487
rect 28859 15453 28871 15487
rect 28994 15484 29000 15496
rect 28955 15456 29000 15484
rect 28813 15447 28871 15453
rect 27062 15416 27068 15428
rect 26160 15388 27068 15416
rect 27062 15376 27068 15388
rect 27120 15376 27126 15428
rect 27522 15416 27528 15428
rect 27483 15388 27528 15416
rect 27522 15376 27528 15388
rect 27580 15376 27586 15428
rect 28552 15416 28580 15444
rect 28828 15416 28856 15447
rect 28994 15444 29000 15456
rect 29052 15444 29058 15496
rect 29089 15487 29147 15493
rect 29089 15453 29101 15487
rect 29135 15453 29147 15487
rect 29089 15447 29147 15453
rect 29917 15487 29975 15493
rect 29917 15453 29929 15487
rect 29963 15484 29975 15487
rect 30190 15484 30196 15496
rect 29963 15456 30196 15484
rect 29963 15453 29975 15456
rect 29917 15447 29975 15453
rect 28552 15388 28856 15416
rect 29104 15416 29132 15447
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 30834 15444 30840 15496
rect 30892 15484 30898 15496
rect 31297 15487 31355 15493
rect 31297 15484 31309 15487
rect 30892 15456 31309 15484
rect 30892 15444 30898 15456
rect 31297 15453 31309 15456
rect 31343 15484 31355 15487
rect 31386 15484 31392 15496
rect 31343 15456 31392 15484
rect 31343 15453 31355 15456
rect 31297 15447 31355 15453
rect 31386 15444 31392 15456
rect 31444 15444 31450 15496
rect 32125 15487 32183 15493
rect 32125 15453 32137 15487
rect 32171 15484 32183 15487
rect 32214 15484 32220 15496
rect 32171 15456 32220 15484
rect 32171 15453 32183 15456
rect 32125 15447 32183 15453
rect 32214 15444 32220 15456
rect 32272 15444 32278 15496
rect 32950 15484 32956 15496
rect 32911 15456 32956 15484
rect 32950 15444 32956 15456
rect 33008 15444 33014 15496
rect 33229 15487 33287 15493
rect 33229 15453 33241 15487
rect 33275 15484 33287 15487
rect 33318 15484 33324 15496
rect 33275 15456 33324 15484
rect 33275 15453 33287 15456
rect 33229 15447 33287 15453
rect 33318 15444 33324 15456
rect 33376 15444 33382 15496
rect 34146 15444 34152 15496
rect 34204 15484 34210 15496
rect 35084 15493 35112 15524
rect 35161 15521 35173 15555
rect 35207 15552 35219 15555
rect 36354 15552 36360 15564
rect 35207 15524 35388 15552
rect 35207 15521 35219 15524
rect 35161 15515 35219 15521
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34204 15456 34897 15484
rect 34204 15444 34210 15456
rect 34885 15453 34897 15456
rect 34931 15453 34943 15487
rect 34885 15447 34943 15453
rect 35069 15487 35127 15493
rect 35069 15453 35081 15487
rect 35115 15453 35127 15487
rect 35069 15447 35127 15453
rect 35253 15487 35311 15493
rect 35253 15453 35265 15487
rect 35299 15453 35311 15487
rect 35253 15447 35311 15453
rect 30926 15416 30932 15428
rect 29104 15388 30932 15416
rect 30926 15376 30932 15388
rect 30984 15376 30990 15428
rect 31018 15376 31024 15428
rect 31076 15416 31082 15428
rect 32306 15416 32312 15428
rect 31076 15388 31169 15416
rect 32267 15388 32312 15416
rect 31076 15376 31082 15388
rect 32306 15376 32312 15388
rect 32364 15376 32370 15428
rect 34790 15376 34796 15428
rect 34848 15416 34854 15428
rect 35268 15416 35296 15447
rect 34848 15388 35296 15416
rect 34848 15376 34854 15388
rect 22281 15351 22339 15357
rect 22281 15317 22293 15351
rect 22327 15348 22339 15351
rect 22370 15348 22376 15360
rect 22327 15320 22376 15348
rect 22327 15317 22339 15320
rect 22281 15311 22339 15317
rect 22370 15308 22376 15320
rect 22428 15308 22434 15360
rect 23290 15308 23296 15360
rect 23348 15348 23354 15360
rect 23385 15351 23443 15357
rect 23385 15348 23397 15351
rect 23348 15320 23397 15348
rect 23348 15308 23354 15320
rect 23385 15317 23397 15320
rect 23431 15317 23443 15351
rect 23385 15311 23443 15317
rect 28537 15351 28595 15357
rect 28537 15317 28549 15351
rect 28583 15348 28595 15351
rect 28626 15348 28632 15360
rect 28583 15320 28632 15348
rect 28583 15317 28595 15320
rect 28537 15311 28595 15317
rect 28626 15308 28632 15320
rect 28684 15308 28690 15360
rect 28902 15308 28908 15360
rect 28960 15348 28966 15360
rect 31036 15348 31064 15376
rect 28960 15320 31064 15348
rect 31205 15351 31263 15357
rect 28960 15308 28966 15320
rect 31205 15317 31217 15351
rect 31251 15348 31263 15351
rect 31294 15348 31300 15360
rect 31251 15320 31300 15348
rect 31251 15317 31263 15320
rect 31205 15311 31263 15317
rect 31294 15308 31300 15320
rect 31352 15308 31358 15360
rect 33137 15351 33195 15357
rect 33137 15317 33149 15351
rect 33183 15348 33195 15351
rect 33410 15348 33416 15360
rect 33183 15320 33416 15348
rect 33183 15317 33195 15320
rect 33137 15311 33195 15317
rect 33410 15308 33416 15320
rect 33468 15308 33474 15360
rect 34330 15348 34336 15360
rect 34291 15320 34336 15348
rect 34330 15308 34336 15320
rect 34388 15308 34394 15360
rect 34698 15308 34704 15360
rect 34756 15348 34762 15360
rect 35360 15348 35388 15524
rect 36280 15524 36360 15552
rect 35437 15487 35495 15493
rect 35437 15453 35449 15487
rect 35483 15453 35495 15487
rect 35437 15447 35495 15453
rect 35452 15416 35480 15447
rect 35894 15444 35900 15496
rect 35952 15484 35958 15496
rect 36280 15493 36308 15524
rect 36354 15512 36360 15524
rect 36412 15512 36418 15564
rect 39022 15552 39028 15564
rect 38983 15524 39028 15552
rect 39022 15512 39028 15524
rect 39080 15512 39086 15564
rect 42981 15555 43039 15561
rect 42981 15521 42993 15555
rect 43027 15552 43039 15555
rect 44836 15552 44864 15580
rect 45370 15552 45376 15564
rect 43027 15524 44864 15552
rect 45331 15524 45376 15552
rect 43027 15521 43039 15524
rect 42981 15515 43039 15521
rect 45370 15512 45376 15524
rect 45428 15512 45434 15564
rect 46106 15552 46112 15564
rect 45480 15524 46112 15552
rect 36265 15487 36323 15493
rect 36265 15484 36277 15487
rect 35952 15456 36277 15484
rect 35952 15444 35958 15456
rect 36265 15453 36277 15456
rect 36311 15453 36323 15487
rect 36630 15484 36636 15496
rect 36591 15456 36636 15484
rect 36265 15447 36323 15453
rect 36630 15444 36636 15456
rect 36688 15444 36694 15496
rect 37185 15487 37243 15493
rect 37185 15453 37197 15487
rect 37231 15484 37243 15487
rect 37645 15487 37703 15493
rect 37645 15484 37657 15487
rect 37231 15456 37657 15484
rect 37231 15453 37243 15456
rect 37185 15447 37243 15453
rect 37645 15453 37657 15456
rect 37691 15484 37703 15487
rect 37826 15484 37832 15496
rect 37691 15456 37832 15484
rect 37691 15453 37703 15456
rect 37645 15447 37703 15453
rect 36354 15416 36360 15428
rect 35452 15388 36360 15416
rect 36354 15376 36360 15388
rect 36412 15376 36418 15428
rect 36446 15376 36452 15428
rect 36504 15416 36510 15428
rect 36504 15388 36549 15416
rect 36504 15376 36510 15388
rect 37200 15348 37228 15447
rect 37826 15444 37832 15456
rect 37884 15444 37890 15496
rect 37921 15487 37979 15493
rect 37921 15453 37933 15487
rect 37967 15484 37979 15487
rect 39114 15484 39120 15496
rect 37967 15456 39120 15484
rect 37967 15453 37979 15456
rect 37921 15447 37979 15453
rect 39114 15444 39120 15456
rect 39172 15444 39178 15496
rect 43165 15487 43223 15493
rect 43165 15453 43177 15487
rect 43211 15453 43223 15487
rect 43165 15447 43223 15453
rect 38654 15376 38660 15428
rect 38712 15416 38718 15428
rect 38933 15419 38991 15425
rect 38933 15416 38945 15419
rect 38712 15388 38945 15416
rect 38712 15376 38718 15388
rect 38933 15385 38945 15388
rect 38979 15416 38991 15419
rect 39942 15416 39948 15428
rect 38979 15388 39948 15416
rect 38979 15385 38991 15388
rect 38933 15379 38991 15385
rect 39942 15376 39948 15388
rect 40000 15376 40006 15428
rect 42518 15376 42524 15428
rect 42576 15416 42582 15428
rect 43180 15416 43208 15447
rect 43254 15444 43260 15496
rect 43312 15484 43318 15496
rect 45189 15487 45247 15493
rect 45189 15484 45201 15487
rect 43312 15456 45201 15484
rect 43312 15444 43318 15456
rect 45189 15453 45201 15456
rect 45235 15453 45247 15487
rect 45189 15447 45247 15453
rect 42576 15388 43208 15416
rect 42576 15376 42582 15388
rect 43622 15376 43628 15428
rect 43680 15416 43686 15428
rect 43993 15419 44051 15425
rect 43993 15416 44005 15419
rect 43680 15388 44005 15416
rect 43680 15376 43686 15388
rect 43993 15385 44005 15388
rect 44039 15416 44051 15419
rect 45480 15416 45508 15524
rect 46106 15512 46112 15524
rect 46164 15512 46170 15564
rect 46308 15552 46336 15592
rect 46477 15623 46535 15629
rect 46477 15589 46489 15623
rect 46523 15620 46535 15623
rect 47946 15620 47952 15632
rect 46523 15592 47952 15620
rect 46523 15589 46535 15592
rect 46477 15583 46535 15589
rect 47946 15580 47952 15592
rect 48004 15580 48010 15632
rect 46216 15524 46336 15552
rect 46385 15555 46443 15561
rect 45557 15487 45615 15493
rect 45557 15453 45569 15487
rect 45603 15453 45615 15487
rect 46216 15484 46244 15524
rect 46385 15521 46397 15555
rect 46431 15552 46443 15555
rect 46658 15552 46664 15564
rect 46431 15524 46664 15552
rect 46431 15521 46443 15524
rect 46385 15515 46443 15521
rect 46658 15512 46664 15524
rect 46716 15512 46722 15564
rect 47394 15552 47400 15564
rect 47355 15524 47400 15552
rect 47394 15512 47400 15524
rect 47452 15512 47458 15564
rect 47486 15512 47492 15564
rect 47544 15552 47550 15564
rect 47673 15555 47731 15561
rect 47544 15524 47589 15552
rect 47544 15512 47550 15524
rect 47673 15521 47685 15555
rect 47719 15552 47731 15555
rect 47762 15552 47768 15564
rect 47719 15524 47768 15552
rect 47719 15521 47731 15524
rect 47673 15515 47731 15521
rect 47762 15512 47768 15524
rect 47820 15512 47826 15564
rect 48286 15552 48314 15660
rect 48682 15648 48688 15700
rect 48740 15688 48746 15700
rect 50154 15688 50160 15700
rect 48740 15660 50160 15688
rect 48740 15648 48746 15660
rect 50154 15648 50160 15660
rect 50212 15648 50218 15700
rect 50614 15648 50620 15700
rect 50672 15688 50678 15700
rect 50801 15691 50859 15697
rect 50801 15688 50813 15691
rect 50672 15660 50813 15688
rect 50672 15648 50678 15660
rect 50801 15657 50813 15660
rect 50847 15657 50859 15691
rect 50801 15651 50859 15657
rect 51626 15648 51632 15700
rect 51684 15688 51690 15700
rect 51905 15691 51963 15697
rect 51905 15688 51917 15691
rect 51684 15660 51917 15688
rect 51684 15648 51690 15660
rect 51905 15657 51917 15660
rect 51951 15657 51963 15691
rect 54938 15688 54944 15700
rect 54899 15660 54944 15688
rect 51905 15651 51963 15657
rect 54938 15648 54944 15660
rect 54996 15648 55002 15700
rect 57514 15688 57520 15700
rect 57475 15660 57520 15688
rect 57514 15648 57520 15660
rect 57572 15648 57578 15700
rect 50062 15580 50068 15632
rect 50120 15620 50126 15632
rect 51810 15620 51816 15632
rect 50120 15592 51816 15620
rect 50120 15580 50126 15592
rect 51810 15580 51816 15592
rect 51868 15620 51874 15632
rect 56778 15620 56784 15632
rect 51868 15592 56784 15620
rect 51868 15580 51874 15592
rect 51261 15555 51319 15561
rect 51261 15552 51273 15555
rect 48286 15524 51273 15552
rect 51261 15521 51273 15524
rect 51307 15552 51319 15555
rect 51902 15552 51908 15564
rect 51307 15524 51908 15552
rect 51307 15521 51319 15524
rect 51261 15515 51319 15521
rect 51902 15512 51908 15524
rect 51960 15512 51966 15564
rect 52380 15561 52408 15592
rect 56778 15580 56784 15592
rect 56836 15580 56842 15632
rect 52365 15555 52423 15561
rect 52365 15521 52377 15555
rect 52411 15521 52423 15555
rect 56594 15552 56600 15564
rect 52365 15515 52423 15521
rect 54128 15524 56600 15552
rect 46293 15487 46351 15493
rect 46293 15484 46305 15487
rect 46216 15456 46305 15484
rect 45557 15447 45615 15453
rect 46293 15453 46305 15456
rect 46339 15453 46351 15487
rect 46293 15447 46351 15453
rect 46569 15487 46627 15493
rect 46569 15453 46581 15487
rect 46615 15484 46627 15487
rect 46842 15484 46848 15496
rect 46615 15456 46848 15484
rect 46615 15453 46627 15456
rect 46569 15447 46627 15453
rect 44039 15388 45508 15416
rect 45572 15416 45600 15447
rect 46842 15444 46848 15456
rect 46900 15484 46906 15496
rect 47026 15484 47032 15496
rect 46900 15456 47032 15484
rect 46900 15444 46906 15456
rect 47026 15444 47032 15456
rect 47084 15444 47090 15496
rect 47578 15484 47584 15496
rect 47539 15456 47584 15484
rect 47578 15444 47584 15456
rect 47636 15444 47642 15496
rect 48222 15444 48228 15496
rect 48280 15484 48286 15496
rect 50341 15487 50399 15493
rect 49252 15484 49464 15486
rect 50341 15484 50353 15487
rect 48280 15458 50353 15484
rect 48280 15456 49280 15458
rect 49436 15456 50353 15458
rect 48280 15444 48286 15456
rect 50341 15453 50353 15456
rect 50387 15453 50399 15487
rect 50341 15447 50399 15453
rect 50617 15487 50675 15493
rect 50617 15453 50629 15487
rect 50663 15484 50675 15487
rect 50706 15484 50712 15496
rect 50663 15456 50712 15484
rect 50663 15453 50675 15456
rect 50617 15447 50675 15453
rect 50706 15444 50712 15456
rect 50764 15444 50770 15496
rect 52089 15487 52147 15493
rect 52089 15453 52101 15487
rect 52135 15453 52147 15487
rect 52270 15484 52276 15496
rect 52231 15456 52276 15484
rect 52089 15447 52147 15453
rect 47394 15416 47400 15428
rect 45572 15388 47400 15416
rect 44039 15385 44051 15388
rect 43993 15379 44051 15385
rect 47394 15376 47400 15388
rect 47452 15376 47458 15428
rect 48317 15419 48375 15425
rect 48317 15416 48329 15419
rect 47504 15388 48329 15416
rect 34756 15320 37228 15348
rect 37829 15351 37887 15357
rect 34756 15308 34762 15320
rect 37829 15317 37841 15351
rect 37875 15348 37887 15351
rect 38746 15348 38752 15360
rect 37875 15320 38752 15348
rect 37875 15317 37887 15320
rect 37829 15311 37887 15317
rect 38746 15308 38752 15320
rect 38804 15308 38810 15360
rect 38841 15351 38899 15357
rect 38841 15317 38853 15351
rect 38887 15348 38899 15351
rect 39390 15348 39396 15360
rect 38887 15320 39396 15348
rect 38887 15317 38899 15320
rect 38841 15311 38899 15317
rect 39390 15308 39396 15320
rect 39448 15348 39454 15360
rect 40037 15351 40095 15357
rect 40037 15348 40049 15351
rect 39448 15320 40049 15348
rect 39448 15308 39454 15320
rect 40037 15317 40049 15320
rect 40083 15348 40095 15351
rect 40862 15348 40868 15360
rect 40083 15320 40868 15348
rect 40083 15317 40095 15320
rect 40037 15311 40095 15317
rect 40862 15308 40868 15320
rect 40920 15308 40926 15360
rect 45278 15348 45284 15360
rect 45239 15320 45284 15348
rect 45278 15308 45284 15320
rect 45336 15308 45342 15360
rect 45465 15351 45523 15357
rect 45465 15317 45477 15351
rect 45511 15348 45523 15351
rect 45646 15348 45652 15360
rect 45511 15320 45652 15348
rect 45511 15317 45523 15320
rect 45465 15311 45523 15317
rect 45646 15308 45652 15320
rect 45704 15308 45710 15360
rect 45738 15308 45744 15360
rect 45796 15348 45802 15360
rect 46198 15348 46204 15360
rect 45796 15320 46204 15348
rect 45796 15308 45802 15320
rect 46198 15308 46204 15320
rect 46256 15308 46262 15360
rect 46750 15308 46756 15360
rect 46808 15348 46814 15360
rect 47504 15348 47532 15388
rect 48317 15385 48329 15388
rect 48363 15416 48375 15419
rect 48869 15419 48927 15425
rect 48869 15416 48881 15419
rect 48363 15388 48881 15416
rect 48363 15385 48375 15388
rect 48317 15379 48375 15385
rect 48869 15385 48881 15388
rect 48915 15385 48927 15419
rect 48869 15379 48927 15385
rect 47854 15348 47860 15360
rect 46808 15320 47532 15348
rect 47815 15320 47860 15348
rect 46808 15308 46814 15320
rect 47854 15308 47860 15320
rect 47912 15308 47918 15360
rect 48884 15348 48912 15379
rect 49234 15376 49240 15428
rect 49292 15416 49298 15428
rect 49421 15419 49479 15425
rect 49421 15416 49433 15419
rect 49292 15388 49433 15416
rect 49292 15376 49298 15388
rect 49421 15385 49433 15388
rect 49467 15385 49479 15419
rect 49421 15379 49479 15385
rect 49605 15419 49663 15425
rect 49605 15385 49617 15419
rect 49651 15416 49663 15419
rect 49970 15416 49976 15428
rect 49651 15388 49976 15416
rect 49651 15385 49663 15388
rect 49605 15379 49663 15385
rect 49970 15376 49976 15388
rect 50028 15376 50034 15428
rect 52104 15416 52132 15447
rect 52270 15444 52276 15456
rect 52328 15444 52334 15496
rect 52454 15444 52460 15496
rect 52512 15484 52518 15496
rect 53009 15487 53067 15493
rect 53009 15484 53021 15487
rect 52512 15456 53021 15484
rect 52512 15444 52518 15456
rect 53009 15453 53021 15456
rect 53055 15453 53067 15487
rect 53190 15484 53196 15496
rect 53151 15456 53196 15484
rect 53009 15447 53067 15453
rect 53190 15444 53196 15456
rect 53248 15444 53254 15496
rect 53285 15487 53343 15493
rect 53285 15453 53297 15487
rect 53331 15484 53343 15487
rect 53466 15484 53472 15496
rect 53331 15456 53472 15484
rect 53331 15453 53343 15456
rect 53285 15447 53343 15453
rect 53466 15444 53472 15456
rect 53524 15444 53530 15496
rect 52914 15416 52920 15428
rect 52104 15388 52920 15416
rect 52914 15376 52920 15388
rect 52972 15376 52978 15428
rect 53208 15416 53236 15444
rect 54128 15416 54156 15524
rect 56594 15512 56600 15524
rect 56652 15552 56658 15564
rect 58069 15555 58127 15561
rect 58069 15552 58081 15555
rect 56652 15524 58081 15552
rect 56652 15512 56658 15524
rect 58069 15521 58081 15524
rect 58115 15521 58127 15555
rect 58069 15515 58127 15521
rect 55214 15444 55220 15496
rect 55272 15484 55278 15496
rect 55953 15487 56011 15493
rect 55953 15484 55965 15487
rect 55272 15456 55965 15484
rect 55272 15444 55278 15456
rect 55953 15453 55965 15456
rect 55999 15484 56011 15487
rect 56686 15484 56692 15496
rect 55999 15456 56692 15484
rect 55999 15453 56011 15456
rect 55953 15447 56011 15453
rect 56686 15444 56692 15456
rect 56744 15484 56750 15496
rect 56965 15487 57023 15493
rect 56965 15484 56977 15487
rect 56744 15456 56977 15484
rect 56744 15444 56750 15456
rect 56965 15453 56977 15456
rect 57011 15453 57023 15487
rect 56965 15447 57023 15453
rect 53208 15388 54156 15416
rect 54478 15376 54484 15428
rect 54536 15416 54542 15428
rect 55585 15419 55643 15425
rect 55585 15416 55597 15419
rect 54536 15388 55597 15416
rect 54536 15376 54542 15388
rect 55585 15385 55597 15388
rect 55631 15416 55643 15419
rect 57146 15416 57152 15428
rect 55631 15388 57152 15416
rect 55631 15385 55643 15388
rect 55585 15379 55643 15385
rect 57146 15376 57152 15388
rect 57204 15376 57210 15428
rect 49510 15348 49516 15360
rect 48884 15320 49516 15348
rect 49510 15308 49516 15320
rect 49568 15308 49574 15360
rect 49789 15351 49847 15357
rect 49789 15317 49801 15351
rect 49835 15348 49847 15351
rect 50433 15351 50491 15357
rect 50433 15348 50445 15351
rect 49835 15320 50445 15348
rect 49835 15317 49847 15320
rect 49789 15311 49847 15317
rect 50433 15317 50445 15320
rect 50479 15317 50491 15351
rect 52822 15348 52828 15360
rect 52783 15320 52828 15348
rect 50433 15311 50491 15317
rect 52822 15308 52828 15320
rect 52880 15308 52886 15360
rect 53650 15308 53656 15360
rect 53708 15348 53714 15360
rect 53745 15351 53803 15357
rect 53745 15348 53757 15351
rect 53708 15320 53757 15348
rect 53708 15308 53714 15320
rect 53745 15317 53757 15320
rect 53791 15317 53803 15351
rect 53745 15311 53803 15317
rect 53834 15308 53840 15360
rect 53892 15348 53898 15360
rect 54297 15351 54355 15357
rect 54297 15348 54309 15351
rect 53892 15320 54309 15348
rect 53892 15308 53898 15320
rect 54297 15317 54309 15320
rect 54343 15317 54355 15351
rect 54297 15311 54355 15317
rect 56226 15308 56232 15360
rect 56284 15348 56290 15360
rect 56413 15351 56471 15357
rect 56413 15348 56425 15351
rect 56284 15320 56425 15348
rect 56284 15308 56290 15320
rect 56413 15317 56425 15320
rect 56459 15317 56471 15351
rect 56413 15311 56471 15317
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 23566 15104 23572 15156
rect 23624 15144 23630 15156
rect 23661 15147 23719 15153
rect 23661 15144 23673 15147
rect 23624 15116 23673 15144
rect 23624 15104 23630 15116
rect 23661 15113 23673 15116
rect 23707 15113 23719 15147
rect 24026 15144 24032 15156
rect 23987 15116 24032 15144
rect 23661 15107 23719 15113
rect 24026 15104 24032 15116
rect 24084 15104 24090 15156
rect 24762 15104 24768 15156
rect 24820 15144 24826 15156
rect 24857 15147 24915 15153
rect 24857 15144 24869 15147
rect 24820 15116 24869 15144
rect 24820 15104 24826 15116
rect 24857 15113 24869 15116
rect 24903 15113 24915 15147
rect 24857 15107 24915 15113
rect 25777 15147 25835 15153
rect 25777 15113 25789 15147
rect 25823 15144 25835 15147
rect 26418 15144 26424 15156
rect 25823 15116 26424 15144
rect 25823 15113 25835 15116
rect 25777 15107 25835 15113
rect 26418 15104 26424 15116
rect 26476 15104 26482 15156
rect 28721 15147 28779 15153
rect 28721 15113 28733 15147
rect 28767 15144 28779 15147
rect 28994 15144 29000 15156
rect 28767 15116 29000 15144
rect 28767 15113 28779 15116
rect 28721 15107 28779 15113
rect 28994 15104 29000 15116
rect 29052 15104 29058 15156
rect 29638 15104 29644 15156
rect 29696 15144 29702 15156
rect 30377 15147 30435 15153
rect 30377 15144 30389 15147
rect 29696 15116 30389 15144
rect 29696 15104 29702 15116
rect 30377 15113 30389 15116
rect 30423 15113 30435 15147
rect 36170 15144 36176 15156
rect 30377 15107 30435 15113
rect 34808 15116 36176 15144
rect 22830 15076 22836 15088
rect 22743 15048 22836 15076
rect 22830 15036 22836 15048
rect 22888 15076 22894 15088
rect 24780 15076 24808 15104
rect 26510 15076 26516 15088
rect 22888 15048 24808 15076
rect 26471 15048 26516 15076
rect 22888 15036 22894 15048
rect 26510 15036 26516 15048
rect 26568 15036 26574 15088
rect 26970 15036 26976 15088
rect 27028 15076 27034 15088
rect 27249 15079 27307 15085
rect 27249 15076 27261 15079
rect 27028 15048 27261 15076
rect 27028 15036 27034 15048
rect 27249 15045 27261 15048
rect 27295 15045 27307 15079
rect 27249 15039 27307 15045
rect 29914 15036 29920 15088
rect 29972 15076 29978 15088
rect 31021 15079 31079 15085
rect 31021 15076 31033 15079
rect 29972 15048 31033 15076
rect 29972 15036 29978 15048
rect 31021 15045 31033 15048
rect 31067 15045 31079 15079
rect 31021 15039 31079 15045
rect 31110 15036 31116 15088
rect 31168 15076 31174 15088
rect 31386 15076 31392 15088
rect 31168 15048 31392 15076
rect 31168 15036 31174 15048
rect 31386 15036 31392 15048
rect 31444 15076 31450 15088
rect 32861 15079 32919 15085
rect 32861 15076 32873 15079
rect 31444 15048 32873 15076
rect 31444 15036 31450 15048
rect 32861 15045 32873 15048
rect 32907 15045 32919 15079
rect 32861 15039 32919 15045
rect 34057 15079 34115 15085
rect 34057 15045 34069 15079
rect 34103 15076 34115 15079
rect 34422 15076 34428 15088
rect 34103 15048 34428 15076
rect 34103 15045 34115 15048
rect 34057 15039 34115 15045
rect 34422 15036 34428 15048
rect 34480 15076 34486 15088
rect 34701 15079 34759 15085
rect 34701 15076 34713 15079
rect 34480 15048 34713 15076
rect 34480 15036 34486 15048
rect 34701 15045 34713 15048
rect 34747 15045 34759 15079
rect 34701 15039 34759 15045
rect 21358 14968 21364 15020
rect 21416 15008 21422 15020
rect 22465 15011 22523 15017
rect 22465 15008 22477 15011
rect 21416 14980 22477 15008
rect 21416 14968 21422 14980
rect 22465 14977 22477 14980
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 25498 14968 25504 15020
rect 25556 15008 25562 15020
rect 25593 15011 25651 15017
rect 25593 15008 25605 15011
rect 25556 14980 25605 15008
rect 25556 14968 25562 14980
rect 25593 14977 25605 14980
rect 25639 15008 25651 15011
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 25639 14980 26249 15008
rect 25639 14977 25651 14980
rect 25593 14971 25651 14977
rect 26237 14977 26249 14980
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 26329 15011 26387 15017
rect 26329 14977 26341 15011
rect 26375 14977 26387 15011
rect 26329 14971 26387 14977
rect 24118 14940 24124 14952
rect 24079 14912 24124 14940
rect 24118 14900 24124 14912
rect 24176 14900 24182 14952
rect 24302 14940 24308 14952
rect 24263 14912 24308 14940
rect 24302 14900 24308 14912
rect 24360 14900 24366 14952
rect 24762 14900 24768 14952
rect 24820 14940 24826 14952
rect 25409 14943 25467 14949
rect 25409 14940 25421 14943
rect 24820 14912 25421 14940
rect 24820 14900 24826 14912
rect 25409 14909 25421 14912
rect 25455 14940 25467 14943
rect 26344 14940 26372 14971
rect 27062 14968 27068 15020
rect 27120 15008 27126 15020
rect 27433 15011 27491 15017
rect 27433 15008 27445 15011
rect 27120 14980 27445 15008
rect 27120 14968 27126 14980
rect 27433 14977 27445 14980
rect 27479 14977 27491 15011
rect 27614 15008 27620 15020
rect 27575 14980 27620 15008
rect 27433 14971 27491 14977
rect 27614 14968 27620 14980
rect 27672 14968 27678 15020
rect 27709 15011 27767 15017
rect 27709 14977 27721 15011
rect 27755 15008 27767 15011
rect 27982 15008 27988 15020
rect 27755 14980 27988 15008
rect 27755 14977 27767 14980
rect 27709 14971 27767 14977
rect 27982 14968 27988 14980
rect 28040 14968 28046 15020
rect 28810 14968 28816 15020
rect 28868 15008 28874 15020
rect 28905 15011 28963 15017
rect 28905 15008 28917 15011
rect 28868 14980 28917 15008
rect 28868 14968 28874 14980
rect 28905 14977 28917 14980
rect 28951 14977 28963 15011
rect 30006 15008 30012 15020
rect 29967 14980 30012 15008
rect 28905 14971 28963 14977
rect 30006 14968 30012 14980
rect 30064 14968 30070 15020
rect 30098 14968 30104 15020
rect 30156 15008 30162 15020
rect 30193 15011 30251 15017
rect 30193 15008 30205 15011
rect 30156 14980 30205 15008
rect 30156 14968 30162 14980
rect 30193 14977 30205 14980
rect 30239 14977 30251 15011
rect 30193 14971 30251 14977
rect 30926 14968 30932 15020
rect 30984 15008 30990 15020
rect 31610 15011 31668 15017
rect 31610 15008 31622 15011
rect 30984 14980 31622 15008
rect 30984 14968 30990 14980
rect 29178 14940 29184 14952
rect 25455 14912 26372 14940
rect 29139 14912 29184 14940
rect 25455 14909 25467 14912
rect 25409 14903 25467 14909
rect 29178 14900 29184 14912
rect 29236 14900 29242 14952
rect 31389 14943 31447 14949
rect 31389 14909 31401 14943
rect 31435 14909 31447 14943
rect 31496 14940 31524 14980
rect 31610 14977 31622 14980
rect 31656 14977 31668 15011
rect 31610 14971 31668 14977
rect 31757 15011 31815 15017
rect 31757 14977 31769 15011
rect 31803 15008 31815 15011
rect 31846 15008 31852 15020
rect 31803 14980 31852 15008
rect 31803 14977 31815 14980
rect 31757 14971 31815 14977
rect 31846 14968 31852 14980
rect 31904 15008 31910 15020
rect 32214 15008 32220 15020
rect 31904 14980 32220 15008
rect 31904 14968 31910 14980
rect 32214 14968 32220 14980
rect 32272 14968 32278 15020
rect 34330 14968 34336 15020
rect 34388 15008 34394 15020
rect 34517 15011 34575 15017
rect 34517 15008 34529 15011
rect 34388 14980 34529 15008
rect 34388 14968 34394 14980
rect 34517 14977 34529 14980
rect 34563 15008 34575 15011
rect 34808 15008 34836 15116
rect 36170 15104 36176 15116
rect 36228 15104 36234 15156
rect 36449 15147 36507 15153
rect 36449 15113 36461 15147
rect 36495 15144 36507 15147
rect 36630 15144 36636 15156
rect 36495 15116 36636 15144
rect 36495 15113 36507 15116
rect 36449 15107 36507 15113
rect 36630 15104 36636 15116
rect 36688 15104 36694 15156
rect 37366 15104 37372 15156
rect 37424 15144 37430 15156
rect 37829 15147 37887 15153
rect 37829 15144 37841 15147
rect 37424 15116 37841 15144
rect 37424 15104 37430 15116
rect 37829 15113 37841 15116
rect 37875 15113 37887 15147
rect 37829 15107 37887 15113
rect 38933 15147 38991 15153
rect 38933 15113 38945 15147
rect 38979 15144 38991 15147
rect 39022 15144 39028 15156
rect 38979 15116 39028 15144
rect 38979 15113 38991 15116
rect 38933 15107 38991 15113
rect 39022 15104 39028 15116
rect 39080 15104 39086 15156
rect 41693 15147 41751 15153
rect 41693 15113 41705 15147
rect 41739 15144 41751 15147
rect 41966 15144 41972 15156
rect 41739 15116 41972 15144
rect 41739 15113 41751 15116
rect 41693 15107 41751 15113
rect 41966 15104 41972 15116
rect 42024 15104 42030 15156
rect 43349 15147 43407 15153
rect 43349 15113 43361 15147
rect 43395 15144 43407 15147
rect 43438 15144 43444 15156
rect 43395 15116 43444 15144
rect 43395 15113 43407 15116
rect 43349 15107 43407 15113
rect 43438 15104 43444 15116
rect 43496 15104 43502 15156
rect 43714 15104 43720 15156
rect 43772 15144 43778 15156
rect 44174 15144 44180 15156
rect 43772 15116 44180 15144
rect 43772 15104 43778 15116
rect 44174 15104 44180 15116
rect 44232 15104 44238 15156
rect 44634 15144 44640 15156
rect 44595 15116 44640 15144
rect 44634 15104 44640 15116
rect 44692 15104 44698 15156
rect 45186 15104 45192 15156
rect 45244 15144 45250 15156
rect 45922 15144 45928 15156
rect 45244 15116 45928 15144
rect 45244 15104 45250 15116
rect 45922 15104 45928 15116
rect 45980 15104 45986 15156
rect 47854 15104 47860 15156
rect 47912 15144 47918 15156
rect 47965 15147 48023 15153
rect 47965 15144 47977 15147
rect 47912 15116 47977 15144
rect 47912 15104 47918 15116
rect 47965 15113 47977 15116
rect 48011 15113 48023 15147
rect 47965 15107 48023 15113
rect 48133 15147 48191 15153
rect 48133 15113 48145 15147
rect 48179 15144 48191 15147
rect 48498 15144 48504 15156
rect 48179 15116 48504 15144
rect 48179 15113 48191 15116
rect 48133 15107 48191 15113
rect 48498 15104 48504 15116
rect 48556 15104 48562 15156
rect 49786 15144 49792 15156
rect 48914 15116 49792 15144
rect 39114 15076 39120 15088
rect 35544 15048 39120 15076
rect 34563 14980 34836 15008
rect 34885 15011 34943 15017
rect 34563 14977 34575 14980
rect 34517 14971 34575 14977
rect 34885 14977 34897 15011
rect 34931 15008 34943 15011
rect 35342 15008 35348 15020
rect 34931 14980 35348 15008
rect 34931 14977 34943 14980
rect 34885 14971 34943 14977
rect 35342 14968 35348 14980
rect 35400 14968 35406 15020
rect 35544 15017 35572 15048
rect 39114 15036 39120 15048
rect 39172 15036 39178 15088
rect 39240 15048 39528 15076
rect 35529 15011 35587 15017
rect 35529 14977 35541 15011
rect 35575 14977 35587 15011
rect 36354 15008 36360 15020
rect 36315 14980 36360 15008
rect 35529 14971 35587 14977
rect 36354 14968 36360 14980
rect 36412 14968 36418 15020
rect 36538 14968 36544 15020
rect 36596 15008 36602 15020
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 36596 14980 37473 15008
rect 36596 14968 36602 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37461 14971 37519 14977
rect 37918 14968 37924 15020
rect 37976 15008 37982 15020
rect 39240 15008 39268 15048
rect 37976 14980 39268 15008
rect 37976 14968 37982 14980
rect 39298 14968 39304 15020
rect 39356 15008 39362 15020
rect 39500 15008 39528 15048
rect 39942 15036 39948 15088
rect 40000 15076 40006 15088
rect 40000 15048 40908 15076
rect 40000 15036 40006 15048
rect 40880 15017 40908 15048
rect 41414 15036 41420 15088
rect 41472 15076 41478 15088
rect 41472 15048 46060 15076
rect 41472 15036 41478 15048
rect 40681 15011 40739 15017
rect 40681 15008 40693 15011
rect 39356 14980 39401 15008
rect 39500 14980 40693 15008
rect 39356 14968 39362 14980
rect 40681 14977 40693 14980
rect 40727 14977 40739 15011
rect 40681 14971 40739 14977
rect 40865 15011 40923 15017
rect 40865 14977 40877 15011
rect 40911 14977 40923 15011
rect 43530 15008 43536 15020
rect 43491 14980 43536 15008
rect 40865 14971 40923 14977
rect 43530 14968 43536 14980
rect 43588 14968 43594 15020
rect 43625 15011 43683 15017
rect 43625 14977 43637 15011
rect 43671 14977 43683 15011
rect 43625 14971 43683 14977
rect 32306 14940 32312 14952
rect 31496 14912 32312 14940
rect 31389 14903 31447 14909
rect 26513 14875 26571 14881
rect 26513 14841 26525 14875
rect 26559 14872 26571 14875
rect 28902 14872 28908 14884
rect 26559 14844 28908 14872
rect 26559 14841 26571 14844
rect 26513 14835 26571 14841
rect 28902 14832 28908 14844
rect 28960 14832 28966 14884
rect 21358 14804 21364 14816
rect 21319 14776 21364 14804
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 27522 14764 27528 14816
rect 27580 14804 27586 14816
rect 28258 14804 28264 14816
rect 27580 14776 28264 14804
rect 27580 14764 27586 14776
rect 28258 14764 28264 14776
rect 28316 14764 28322 14816
rect 29089 14807 29147 14813
rect 29089 14773 29101 14807
rect 29135 14804 29147 14807
rect 30190 14804 30196 14816
rect 29135 14776 30196 14804
rect 29135 14773 29147 14776
rect 29089 14767 29147 14773
rect 30190 14764 30196 14776
rect 30248 14764 30254 14816
rect 31404 14804 31432 14903
rect 32306 14900 32312 14912
rect 32364 14900 32370 14952
rect 32401 14943 32459 14949
rect 32401 14909 32413 14943
rect 32447 14940 32459 14943
rect 32674 14940 32680 14952
rect 32447 14912 32680 14940
rect 32447 14909 32459 14912
rect 32401 14903 32459 14909
rect 32674 14900 32680 14912
rect 32732 14940 32738 14952
rect 35618 14940 35624 14952
rect 32732 14912 35624 14940
rect 32732 14900 32738 14912
rect 35618 14900 35624 14912
rect 35676 14940 35682 14952
rect 37553 14943 37611 14949
rect 35676 14912 35940 14940
rect 35676 14900 35682 14912
rect 31481 14875 31539 14881
rect 31481 14841 31493 14875
rect 31527 14872 31539 14875
rect 32490 14872 32496 14884
rect 31527 14844 32496 14872
rect 31527 14841 31539 14844
rect 31481 14835 31539 14841
rect 32490 14832 32496 14844
rect 32548 14832 32554 14884
rect 32582 14832 32588 14884
rect 32640 14872 32646 14884
rect 35437 14875 35495 14881
rect 35437 14872 35449 14875
rect 32640 14844 35449 14872
rect 32640 14832 32646 14844
rect 35437 14841 35449 14844
rect 35483 14872 35495 14875
rect 35802 14872 35808 14884
rect 35483 14844 35808 14872
rect 35483 14841 35495 14844
rect 35437 14835 35495 14841
rect 35802 14832 35808 14844
rect 35860 14832 35866 14884
rect 35912 14872 35940 14912
rect 37553 14909 37565 14943
rect 37599 14940 37611 14943
rect 37734 14940 37740 14952
rect 37599 14912 37740 14940
rect 37599 14909 37611 14912
rect 37553 14903 37611 14909
rect 37734 14900 37740 14912
rect 37792 14940 37798 14952
rect 38286 14940 38292 14952
rect 37792 14912 38292 14940
rect 37792 14900 37798 14912
rect 38286 14900 38292 14912
rect 38344 14900 38350 14952
rect 39114 14940 39120 14952
rect 39075 14912 39120 14940
rect 39114 14900 39120 14912
rect 39172 14900 39178 14952
rect 39209 14943 39267 14949
rect 39209 14909 39221 14943
rect 39255 14909 39267 14943
rect 39209 14903 39267 14909
rect 39393 14943 39451 14949
rect 39393 14909 39405 14943
rect 39439 14940 39451 14943
rect 39482 14940 39488 14952
rect 39439 14912 39488 14940
rect 39439 14909 39451 14912
rect 39393 14903 39451 14909
rect 35912 14844 38654 14872
rect 31754 14804 31760 14816
rect 31404 14776 31760 14804
rect 31754 14764 31760 14776
rect 31812 14764 31818 14816
rect 32858 14764 32864 14816
rect 32916 14804 32922 14816
rect 33413 14807 33471 14813
rect 33413 14804 33425 14807
rect 32916 14776 33425 14804
rect 32916 14764 32922 14776
rect 33413 14773 33425 14776
rect 33459 14804 33471 14807
rect 34698 14804 34704 14816
rect 33459 14776 34704 14804
rect 33459 14773 33471 14776
rect 33413 14767 33471 14773
rect 34698 14764 34704 14776
rect 34756 14764 34762 14816
rect 37458 14804 37464 14816
rect 37419 14776 37464 14804
rect 37458 14764 37464 14776
rect 37516 14764 37522 14816
rect 38194 14764 38200 14816
rect 38252 14804 38258 14816
rect 38289 14807 38347 14813
rect 38289 14804 38301 14807
rect 38252 14776 38301 14804
rect 38252 14764 38258 14776
rect 38289 14773 38301 14776
rect 38335 14773 38347 14807
rect 38626 14804 38654 14844
rect 38838 14832 38844 14884
rect 38896 14872 38902 14884
rect 39224 14872 39252 14903
rect 39482 14900 39488 14912
rect 39540 14900 39546 14952
rect 43640 14940 43668 14971
rect 43714 14968 43720 15020
rect 43772 15008 43778 15020
rect 44818 15008 44824 15020
rect 43772 14980 43817 15008
rect 44779 14980 44824 15008
rect 43772 14968 43778 14980
rect 44818 14968 44824 14980
rect 44876 14968 44882 15020
rect 44910 14968 44916 15020
rect 44968 15008 44974 15020
rect 45097 15011 45155 15017
rect 44968 14980 45013 15008
rect 44968 14968 44974 14980
rect 45097 14977 45109 15011
rect 45143 15008 45155 15011
rect 45186 15008 45192 15020
rect 45143 14980 45192 15008
rect 45143 14977 45155 14980
rect 45097 14971 45155 14977
rect 45186 14968 45192 14980
rect 45244 14968 45250 15020
rect 45646 15008 45652 15020
rect 45607 14980 45652 15008
rect 45646 14968 45652 14980
rect 45704 14968 45710 15020
rect 45738 14968 45744 15020
rect 45796 15008 45802 15020
rect 45922 15008 45928 15020
rect 45796 14980 45841 15008
rect 45883 14980 45928 15008
rect 45796 14968 45802 14980
rect 45922 14968 45928 14980
rect 45980 14968 45986 15020
rect 46032 15017 46060 15048
rect 46198 15036 46204 15088
rect 46256 15076 46262 15088
rect 46937 15079 46995 15085
rect 46937 15076 46949 15079
rect 46256 15048 46949 15076
rect 46256 15036 46262 15048
rect 46937 15045 46949 15048
rect 46983 15045 46995 15079
rect 46937 15039 46995 15045
rect 46017 15011 46075 15017
rect 46017 14977 46029 15011
rect 46063 14977 46075 15011
rect 46017 14971 46075 14977
rect 46106 14968 46112 15020
rect 46164 15008 46170 15020
rect 46753 15011 46811 15017
rect 46753 15008 46765 15011
rect 46164 14980 46765 15008
rect 46164 14968 46170 14980
rect 46753 14977 46765 14980
rect 46799 14977 46811 15011
rect 46952 15008 46980 15039
rect 47394 15036 47400 15088
rect 47452 15076 47458 15088
rect 47762 15076 47768 15088
rect 47452 15048 47768 15076
rect 47452 15036 47458 15048
rect 47762 15036 47768 15048
rect 47820 15036 47826 15088
rect 48914 15076 48942 15116
rect 49786 15104 49792 15116
rect 49844 15104 49850 15156
rect 49970 15144 49976 15156
rect 49883 15116 49976 15144
rect 47872 15048 48942 15076
rect 48972 15048 49740 15076
rect 47872 15008 47900 15048
rect 46952 14980 47900 15008
rect 46753 14971 46811 14977
rect 48038 14968 48044 15020
rect 48096 15008 48102 15020
rect 48593 15011 48651 15017
rect 48593 15008 48605 15011
rect 48096 14980 48605 15008
rect 48096 14968 48102 14980
rect 48593 14977 48605 14980
rect 48639 14977 48651 15011
rect 48774 15008 48780 15020
rect 48735 14980 48780 15008
rect 48593 14971 48651 14977
rect 48774 14968 48780 14980
rect 48832 14968 48838 15020
rect 48972 15017 49000 15048
rect 48961 15011 49019 15017
rect 48961 14977 48973 15011
rect 49007 14977 49019 15011
rect 48961 14971 49019 14977
rect 49053 15011 49111 15017
rect 49053 14977 49065 15011
rect 49099 14977 49111 15011
rect 49053 14971 49111 14977
rect 43640 14912 44496 14940
rect 43898 14872 43904 14884
rect 38896 14844 39252 14872
rect 43859 14844 43904 14872
rect 38896 14832 38902 14844
rect 43898 14832 43904 14844
rect 43956 14832 43962 14884
rect 39206 14804 39212 14816
rect 38626 14776 39212 14804
rect 38289 14767 38347 14773
rect 39206 14764 39212 14776
rect 39264 14804 39270 14816
rect 39945 14807 40003 14813
rect 39945 14804 39957 14807
rect 39264 14776 39957 14804
rect 39264 14764 39270 14776
rect 39945 14773 39957 14776
rect 39991 14773 40003 14807
rect 39945 14767 40003 14773
rect 42889 14807 42947 14813
rect 42889 14773 42901 14807
rect 42935 14804 42947 14807
rect 43806 14804 43812 14816
rect 42935 14776 43812 14804
rect 42935 14773 42947 14776
rect 42889 14767 42947 14773
rect 43806 14764 43812 14776
rect 43864 14764 43870 14816
rect 44468 14804 44496 14912
rect 44542 14900 44548 14952
rect 44600 14940 44606 14952
rect 46201 14943 46259 14949
rect 46201 14940 46213 14943
rect 44600 14912 46213 14940
rect 44600 14900 44606 14912
rect 46201 14909 46213 14912
rect 46247 14909 46259 14943
rect 46201 14903 46259 14909
rect 46658 14900 46664 14952
rect 46716 14940 46722 14952
rect 48682 14940 48688 14952
rect 46716 14912 48688 14940
rect 46716 14900 46722 14912
rect 48682 14900 48688 14912
rect 48740 14900 48746 14952
rect 48866 14940 48872 14952
rect 48827 14912 48872 14940
rect 48866 14900 48872 14912
rect 48924 14900 48930 14952
rect 45005 14875 45063 14881
rect 45005 14841 45017 14875
rect 45051 14872 45063 14875
rect 45462 14872 45468 14884
rect 45051 14844 45468 14872
rect 45051 14841 45063 14844
rect 45005 14835 45063 14841
rect 45462 14832 45468 14844
rect 45520 14832 45526 14884
rect 45554 14832 45560 14884
rect 45612 14872 45618 14884
rect 48406 14872 48412 14884
rect 45612 14844 48412 14872
rect 45612 14832 45618 14844
rect 48406 14832 48412 14844
rect 48464 14832 48470 14884
rect 48498 14832 48504 14884
rect 48556 14872 48562 14884
rect 49068 14872 49096 14971
rect 49326 14968 49332 15020
rect 49384 15008 49390 15020
rect 49384 14980 49648 15008
rect 49384 14968 49390 14980
rect 49252 14912 49372 14940
rect 49252 14881 49280 14912
rect 49344 14884 49372 14912
rect 48556 14844 49096 14872
rect 49237 14875 49295 14881
rect 48556 14832 48562 14844
rect 49237 14841 49249 14875
rect 49283 14841 49295 14875
rect 49237 14835 49295 14841
rect 49326 14832 49332 14884
rect 49384 14832 49390 14884
rect 49620 14872 49648 14980
rect 49712 14949 49740 15048
rect 49896 15017 49924 15116
rect 49970 15104 49976 15116
rect 50028 15144 50034 15156
rect 51442 15144 51448 15156
rect 50028 15116 51448 15144
rect 50028 15104 50034 15116
rect 51442 15104 51448 15116
rect 51500 15104 51506 15156
rect 53117 15147 53175 15153
rect 53117 15144 53129 15147
rect 52104 15116 53129 15144
rect 51169 15079 51227 15085
rect 51169 15045 51181 15079
rect 51215 15076 51227 15079
rect 51258 15076 51264 15088
rect 51215 15048 51264 15076
rect 51215 15045 51227 15048
rect 51169 15039 51227 15045
rect 51258 15036 51264 15048
rect 51316 15036 51322 15088
rect 50246 15017 50252 15020
rect 49881 15011 49939 15017
rect 49881 14977 49893 15011
rect 49927 14977 49939 15011
rect 50202 15011 50252 15017
rect 50202 15008 50214 15011
rect 50194 14978 50214 15008
rect 49881 14971 49939 14977
rect 50202 14977 50214 14978
rect 50248 14977 50252 15011
rect 50202 14971 50252 14977
rect 50246 14968 50252 14971
rect 50304 14968 50310 15020
rect 50338 14968 50344 15020
rect 50396 15008 50402 15020
rect 50890 15008 50896 15020
rect 50396 14980 50785 15008
rect 50851 14980 50896 15008
rect 50396 14968 50402 14980
rect 49697 14943 49755 14949
rect 49697 14909 49709 14943
rect 49743 14909 49755 14943
rect 49697 14903 49755 14909
rect 49973 14943 50031 14949
rect 49973 14909 49985 14943
rect 50019 14909 50031 14943
rect 49973 14903 50031 14909
rect 49988 14872 50016 14903
rect 50062 14900 50068 14952
rect 50120 14940 50126 14952
rect 50757 14940 50785 14980
rect 50890 14968 50896 14980
rect 50948 14968 50954 15020
rect 51077 15011 51135 15017
rect 51077 14977 51089 15011
rect 51123 15008 51135 15011
rect 51442 15008 51448 15020
rect 51123 14980 51448 15008
rect 51123 14977 51135 14980
rect 51077 14971 51135 14977
rect 51442 14968 51448 14980
rect 51500 14968 51506 15020
rect 51718 14968 51724 15020
rect 51776 15008 51782 15020
rect 52104 15017 52132 15116
rect 53117 15113 53129 15116
rect 53163 15113 53175 15147
rect 53282 15144 53288 15156
rect 53243 15116 53288 15144
rect 53117 15107 53175 15113
rect 53282 15104 53288 15116
rect 53340 15104 53346 15156
rect 53837 15147 53895 15153
rect 53837 15113 53849 15147
rect 53883 15144 53895 15147
rect 54570 15144 54576 15156
rect 53883 15116 54576 15144
rect 53883 15113 53895 15116
rect 53837 15107 53895 15113
rect 54570 15104 54576 15116
rect 54628 15104 54634 15156
rect 52365 15079 52423 15085
rect 52365 15045 52377 15079
rect 52411 15076 52423 15079
rect 52822 15076 52828 15088
rect 52411 15048 52828 15076
rect 52411 15045 52423 15048
rect 52365 15039 52423 15045
rect 52822 15036 52828 15048
rect 52880 15036 52886 15088
rect 52917 15079 52975 15085
rect 52917 15045 52929 15079
rect 52963 15076 52975 15079
rect 53006 15076 53012 15088
rect 52963 15048 53012 15076
rect 52963 15045 52975 15048
rect 52917 15039 52975 15045
rect 53006 15036 53012 15048
rect 53064 15036 53070 15088
rect 54662 15036 54668 15088
rect 54720 15076 54726 15088
rect 54720 15048 56640 15076
rect 54720 15036 54726 15048
rect 52089 15011 52147 15017
rect 52089 15008 52101 15011
rect 51776 14980 52101 15008
rect 51776 14968 51782 14980
rect 52089 14977 52101 14980
rect 52135 14977 52147 15011
rect 52089 14971 52147 14977
rect 52181 15011 52239 15017
rect 52181 14977 52193 15011
rect 52227 14977 52239 15011
rect 54018 15008 54024 15020
rect 53979 14980 54024 15008
rect 52181 14971 52239 14977
rect 51626 14940 51632 14952
rect 50120 14912 50165 14940
rect 50757 14912 51632 14940
rect 50120 14900 50126 14912
rect 51626 14900 51632 14912
rect 51684 14900 51690 14952
rect 49620 14844 50016 14872
rect 45922 14804 45928 14816
rect 44468 14776 45928 14804
rect 45922 14764 45928 14776
rect 45980 14764 45986 14816
rect 47026 14764 47032 14816
rect 47084 14804 47090 14816
rect 47121 14807 47179 14813
rect 47121 14804 47133 14807
rect 47084 14776 47133 14804
rect 47084 14764 47090 14776
rect 47121 14773 47133 14776
rect 47167 14773 47179 14807
rect 47121 14767 47179 14773
rect 47210 14764 47216 14816
rect 47268 14804 47274 14816
rect 47949 14807 48007 14813
rect 47949 14804 47961 14807
rect 47268 14776 47961 14804
rect 47268 14764 47274 14776
rect 47949 14773 47961 14776
rect 47995 14804 48007 14807
rect 48222 14804 48228 14816
rect 47995 14776 48228 14804
rect 47995 14773 48007 14776
rect 47949 14767 48007 14773
rect 48222 14764 48228 14776
rect 48280 14764 48286 14816
rect 50614 14764 50620 14816
rect 50672 14804 50678 14816
rect 51074 14804 51080 14816
rect 50672 14776 51080 14804
rect 50672 14764 50678 14776
rect 51074 14764 51080 14776
rect 51132 14804 51138 14816
rect 52196 14804 52224 14971
rect 54018 14968 54024 14980
rect 54076 14968 54082 15020
rect 54113 15011 54171 15017
rect 54113 14977 54125 15011
rect 54159 14977 54171 15011
rect 54113 14971 54171 14977
rect 53282 14900 53288 14952
rect 53340 14940 53346 14952
rect 54128 14940 54156 14971
rect 54202 14968 54208 15020
rect 54260 15008 54266 15020
rect 54297 15011 54355 15017
rect 54297 15008 54309 15011
rect 54260 14980 54309 15008
rect 54260 14968 54266 14980
rect 54297 14977 54309 14980
rect 54343 14977 54355 15011
rect 54297 14971 54355 14977
rect 54386 14968 54392 15020
rect 54444 15008 54450 15020
rect 55214 15008 55220 15020
rect 54444 14980 54489 15008
rect 55175 14980 55220 15008
rect 54444 14968 54450 14980
rect 55214 14968 55220 14980
rect 55272 14968 55278 15020
rect 55490 15008 55496 15020
rect 55451 14980 55496 15008
rect 55490 14968 55496 14980
rect 55548 14968 55554 15020
rect 55582 14968 55588 15020
rect 55640 15008 55646 15020
rect 55677 15011 55735 15017
rect 55677 15008 55689 15011
rect 55640 14980 55689 15008
rect 55640 14968 55646 14980
rect 55677 14977 55689 14980
rect 55723 14977 55735 15011
rect 55677 14971 55735 14977
rect 55950 14968 55956 15020
rect 56008 15008 56014 15020
rect 56612 15017 56640 15048
rect 56045 15011 56103 15017
rect 56045 15008 56057 15011
rect 56008 14980 56057 15008
rect 56008 14968 56014 14980
rect 56045 14977 56057 14980
rect 56091 14977 56103 15011
rect 56045 14971 56103 14977
rect 56597 15011 56655 15017
rect 56597 14977 56609 15011
rect 56643 14977 56655 15011
rect 56962 15008 56968 15020
rect 56923 14980 56968 15008
rect 56597 14971 56655 14977
rect 56962 14968 56968 14980
rect 57020 14968 57026 15020
rect 53340 14912 55720 14940
rect 53340 14900 53346 14912
rect 55692 14884 55720 14912
rect 52270 14832 52276 14884
rect 52328 14872 52334 14884
rect 52365 14875 52423 14881
rect 52365 14872 52377 14875
rect 52328 14844 52377 14872
rect 52328 14832 52334 14844
rect 52365 14841 52377 14844
rect 52411 14841 52423 14875
rect 52365 14835 52423 14841
rect 53466 14832 53472 14884
rect 53524 14872 53530 14884
rect 54110 14872 54116 14884
rect 53524 14844 54116 14872
rect 53524 14832 53530 14844
rect 54110 14832 54116 14844
rect 54168 14832 54174 14884
rect 55674 14832 55680 14884
rect 55732 14832 55738 14884
rect 53101 14807 53159 14813
rect 53101 14804 53113 14807
rect 51132 14776 53113 14804
rect 51132 14764 51138 14776
rect 53101 14773 53113 14776
rect 53147 14773 53159 14807
rect 53101 14767 53159 14773
rect 57882 14764 57888 14816
rect 57940 14804 57946 14816
rect 58069 14807 58127 14813
rect 58069 14804 58081 14807
rect 57940 14776 58081 14804
rect 57940 14764 57946 14776
rect 58069 14773 58081 14776
rect 58115 14773 58127 14807
rect 58069 14767 58127 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 24118 14560 24124 14612
rect 24176 14600 24182 14612
rect 24581 14603 24639 14609
rect 24581 14600 24593 14603
rect 24176 14572 24593 14600
rect 24176 14560 24182 14572
rect 24581 14569 24593 14572
rect 24627 14569 24639 14603
rect 24581 14563 24639 14569
rect 26234 14560 26240 14612
rect 26292 14600 26298 14612
rect 26789 14603 26847 14609
rect 26789 14600 26801 14603
rect 26292 14572 26801 14600
rect 26292 14560 26298 14572
rect 26789 14569 26801 14572
rect 26835 14600 26847 14603
rect 27614 14600 27620 14612
rect 26835 14572 27620 14600
rect 26835 14569 26847 14572
rect 26789 14563 26847 14569
rect 27614 14560 27620 14572
rect 27672 14600 27678 14612
rect 28534 14600 28540 14612
rect 27672 14572 28540 14600
rect 27672 14560 27678 14572
rect 28534 14560 28540 14572
rect 28592 14600 28598 14612
rect 29914 14600 29920 14612
rect 28592 14572 29920 14600
rect 28592 14560 28598 14572
rect 29914 14560 29920 14572
rect 29972 14560 29978 14612
rect 31849 14603 31907 14609
rect 31849 14569 31861 14603
rect 31895 14600 31907 14603
rect 32306 14600 32312 14612
rect 31895 14572 32312 14600
rect 31895 14569 31907 14572
rect 31849 14563 31907 14569
rect 32306 14560 32312 14572
rect 32364 14560 32370 14612
rect 32398 14560 32404 14612
rect 32456 14600 32462 14612
rect 32953 14603 33011 14609
rect 32953 14600 32965 14603
rect 32456 14572 32965 14600
rect 32456 14560 32462 14572
rect 32953 14569 32965 14572
rect 32999 14569 33011 14603
rect 33410 14600 33416 14612
rect 33371 14572 33416 14600
rect 32953 14563 33011 14569
rect 33410 14560 33416 14572
rect 33468 14560 33474 14612
rect 35434 14560 35440 14612
rect 35492 14600 35498 14612
rect 35529 14603 35587 14609
rect 35529 14600 35541 14603
rect 35492 14572 35541 14600
rect 35492 14560 35498 14572
rect 35529 14569 35541 14572
rect 35575 14569 35587 14603
rect 36538 14600 36544 14612
rect 36499 14572 36544 14600
rect 35529 14563 35587 14569
rect 36538 14560 36544 14572
rect 36596 14560 36602 14612
rect 36725 14603 36783 14609
rect 36725 14569 36737 14603
rect 36771 14569 36783 14603
rect 37918 14600 37924 14612
rect 37879 14572 37924 14600
rect 36725 14563 36783 14569
rect 22557 14535 22615 14541
rect 22557 14501 22569 14535
rect 22603 14532 22615 14535
rect 29086 14532 29092 14544
rect 22603 14504 23060 14532
rect 22603 14501 22615 14504
rect 22557 14495 22615 14501
rect 23032 14473 23060 14504
rect 26344 14504 29092 14532
rect 23017 14467 23075 14473
rect 23017 14433 23029 14467
rect 23063 14433 23075 14467
rect 23017 14427 23075 14433
rect 25133 14467 25191 14473
rect 25133 14433 25145 14467
rect 25179 14433 25191 14467
rect 25133 14427 25191 14433
rect 22370 14396 22376 14408
rect 22331 14368 22376 14396
rect 22370 14356 22376 14368
rect 22428 14356 22434 14408
rect 23290 14396 23296 14408
rect 23251 14368 23296 14396
rect 23290 14356 23296 14368
rect 23348 14356 23354 14408
rect 24670 14356 24676 14408
rect 24728 14396 24734 14408
rect 25148 14396 25176 14427
rect 24728 14368 25176 14396
rect 24728 14356 24734 14368
rect 24946 14328 24952 14340
rect 24907 14300 24952 14328
rect 24946 14288 24952 14300
rect 25004 14288 25010 14340
rect 26344 14328 26372 14504
rect 29086 14492 29092 14504
rect 29144 14492 29150 14544
rect 32674 14492 32680 14544
rect 32732 14492 32738 14544
rect 32951 14504 34099 14532
rect 27341 14467 27399 14473
rect 27341 14433 27353 14467
rect 27387 14464 27399 14467
rect 27706 14464 27712 14476
rect 27387 14436 27712 14464
rect 27387 14433 27399 14436
rect 27341 14427 27399 14433
rect 27706 14424 27712 14436
rect 27764 14464 27770 14476
rect 28166 14464 28172 14476
rect 27764 14436 28172 14464
rect 27764 14424 27770 14436
rect 28166 14424 28172 14436
rect 28224 14424 28230 14476
rect 28258 14424 28264 14476
rect 28316 14464 28322 14476
rect 28353 14467 28411 14473
rect 28353 14464 28365 14467
rect 28316 14436 28365 14464
rect 28316 14424 28322 14436
rect 28353 14433 28365 14436
rect 28399 14464 28411 14467
rect 32692 14464 32720 14492
rect 28399 14436 31156 14464
rect 28399 14433 28411 14436
rect 28353 14427 28411 14433
rect 31128 14408 31156 14436
rect 31496 14436 32720 14464
rect 27525 14399 27583 14405
rect 27525 14365 27537 14399
rect 27571 14365 27583 14399
rect 27525 14359 27583 14365
rect 26510 14328 26516 14340
rect 25056 14300 26372 14328
rect 26471 14300 26516 14328
rect 25056 14269 25084 14300
rect 26510 14288 26516 14300
rect 26568 14328 26574 14340
rect 27540 14328 27568 14359
rect 27614 14356 27620 14408
rect 27672 14396 27678 14408
rect 27801 14399 27859 14405
rect 27801 14396 27813 14399
rect 27672 14368 27813 14396
rect 27672 14356 27678 14368
rect 27801 14365 27813 14368
rect 27847 14365 27859 14399
rect 27801 14359 27859 14365
rect 31110 14356 31116 14408
rect 31168 14396 31174 14408
rect 31205 14399 31263 14405
rect 31205 14396 31217 14399
rect 31168 14368 31217 14396
rect 31168 14356 31174 14368
rect 31205 14365 31217 14368
rect 31251 14365 31263 14399
rect 31386 14396 31392 14408
rect 31347 14368 31392 14396
rect 31205 14359 31263 14365
rect 31386 14356 31392 14368
rect 31444 14356 31450 14408
rect 31496 14405 31524 14436
rect 31481 14399 31539 14405
rect 31481 14365 31493 14399
rect 31527 14365 31539 14399
rect 31481 14359 31539 14365
rect 31570 14356 31576 14408
rect 31628 14396 31634 14408
rect 32306 14396 32312 14408
rect 31628 14368 31673 14396
rect 32267 14368 32312 14396
rect 31628 14356 31634 14368
rect 32306 14356 32312 14368
rect 32364 14356 32370 14408
rect 32490 14396 32496 14408
rect 32451 14368 32496 14396
rect 32490 14356 32496 14368
rect 32548 14356 32554 14408
rect 32582 14356 32588 14408
rect 32640 14396 32646 14408
rect 32723 14399 32781 14405
rect 32640 14368 32685 14396
rect 32640 14356 32646 14368
rect 32723 14365 32735 14399
rect 32769 14396 32781 14399
rect 32858 14396 32864 14408
rect 32769 14368 32864 14396
rect 32769 14365 32781 14368
rect 32723 14359 32781 14365
rect 32858 14356 32864 14368
rect 32916 14356 32922 14408
rect 26568 14300 27568 14328
rect 27709 14331 27767 14337
rect 26568 14288 26574 14300
rect 27709 14297 27721 14331
rect 27755 14328 27767 14331
rect 28258 14328 28264 14340
rect 27755 14300 28264 14328
rect 27755 14297 27767 14300
rect 27709 14291 27767 14297
rect 24029 14263 24087 14269
rect 24029 14229 24041 14263
rect 24075 14260 24087 14263
rect 25041 14263 25099 14269
rect 25041 14260 25053 14263
rect 24075 14232 25053 14260
rect 24075 14229 24087 14232
rect 24029 14223 24087 14229
rect 25041 14229 25053 14232
rect 25087 14229 25099 14263
rect 25041 14223 25099 14229
rect 25961 14263 26019 14269
rect 25961 14229 25973 14263
rect 26007 14260 26019 14263
rect 26142 14260 26148 14272
rect 26007 14232 26148 14260
rect 26007 14229 26019 14232
rect 25961 14223 26019 14229
rect 26142 14220 26148 14232
rect 26200 14260 26206 14272
rect 27724 14260 27752 14291
rect 28258 14288 28264 14300
rect 28316 14288 28322 14340
rect 29546 14328 29552 14340
rect 28368 14300 29552 14328
rect 26200 14232 27752 14260
rect 26200 14220 26206 14232
rect 27890 14220 27896 14272
rect 27948 14260 27954 14272
rect 28368 14260 28396 14300
rect 29546 14288 29552 14300
rect 29604 14328 29610 14340
rect 32951 14328 32979 14504
rect 33778 14424 33784 14476
rect 33836 14424 33842 14476
rect 34071 14464 34099 14504
rect 36262 14492 36268 14544
rect 36320 14532 36326 14544
rect 36740 14532 36768 14563
rect 37918 14560 37924 14572
rect 37976 14560 37982 14612
rect 38378 14600 38384 14612
rect 38339 14572 38384 14600
rect 38378 14560 38384 14572
rect 38436 14560 38442 14612
rect 40586 14600 40592 14612
rect 40547 14572 40592 14600
rect 40586 14560 40592 14572
rect 40644 14560 40650 14612
rect 41414 14560 41420 14612
rect 41472 14600 41478 14612
rect 43070 14600 43076 14612
rect 41472 14572 41517 14600
rect 41892 14572 43076 14600
rect 41472 14560 41478 14572
rect 36320 14504 36768 14532
rect 36320 14492 36326 14504
rect 36814 14492 36820 14544
rect 36872 14532 36878 14544
rect 39482 14532 39488 14544
rect 36872 14504 39488 14532
rect 36872 14492 36878 14504
rect 39482 14492 39488 14504
rect 39540 14492 39546 14544
rect 35342 14464 35348 14476
rect 34071 14436 35112 14464
rect 33689 14399 33747 14405
rect 33600 14377 33658 14383
rect 33600 14343 33612 14377
rect 33646 14343 33658 14377
rect 33689 14365 33701 14399
rect 33735 14393 33747 14399
rect 33796 14393 33824 14424
rect 33735 14365 33824 14393
rect 33885 14399 33943 14405
rect 33885 14365 33897 14399
rect 33931 14365 33943 14399
rect 33689 14359 33747 14365
rect 33885 14359 33943 14365
rect 33975 14399 34033 14405
rect 33975 14365 33987 14399
rect 34021 14396 34033 14399
rect 34071 14396 34099 14436
rect 34882 14396 34888 14408
rect 34021 14368 34099 14396
rect 34843 14368 34888 14396
rect 34021 14365 34033 14368
rect 33975 14359 34033 14365
rect 33600 14340 33658 14343
rect 29604 14300 32979 14328
rect 29604 14288 29610 14300
rect 33594 14288 33600 14340
rect 33652 14288 33658 14340
rect 33888 14272 33916 14359
rect 34882 14356 34888 14368
rect 34940 14356 34946 14408
rect 35084 14405 35112 14436
rect 35176 14436 35348 14464
rect 35176 14405 35204 14436
rect 35342 14424 35348 14436
rect 35400 14424 35406 14476
rect 36354 14424 36360 14476
rect 36412 14464 36418 14476
rect 37461 14467 37519 14473
rect 37461 14464 37473 14467
rect 36412 14436 37473 14464
rect 36412 14424 36418 14436
rect 37461 14433 37473 14436
rect 37507 14464 37519 14467
rect 39298 14464 39304 14476
rect 37507 14436 39304 14464
rect 37507 14433 37519 14436
rect 37461 14427 37519 14433
rect 39298 14424 39304 14436
rect 39356 14424 39362 14476
rect 40405 14467 40463 14473
rect 40405 14433 40417 14467
rect 40451 14464 40463 14467
rect 40586 14464 40592 14476
rect 40451 14436 40592 14464
rect 40451 14433 40463 14436
rect 40405 14427 40463 14433
rect 40586 14424 40592 14436
rect 40644 14424 40650 14476
rect 35069 14399 35127 14405
rect 35069 14365 35081 14399
rect 35115 14365 35127 14399
rect 35069 14359 35127 14365
rect 35161 14399 35219 14405
rect 35161 14365 35173 14399
rect 35207 14365 35219 14399
rect 35161 14359 35219 14365
rect 35253 14399 35311 14405
rect 35253 14365 35265 14399
rect 35299 14396 35311 14399
rect 36372 14396 36400 14424
rect 35299 14368 36400 14396
rect 35299 14365 35311 14368
rect 35253 14359 35311 14365
rect 37550 14356 37556 14408
rect 37608 14396 37614 14408
rect 37737 14399 37795 14405
rect 37608 14368 37653 14396
rect 37608 14356 37614 14368
rect 37737 14365 37749 14399
rect 37783 14365 37795 14399
rect 37737 14359 37795 14365
rect 36081 14331 36139 14337
rect 36081 14297 36093 14331
rect 36127 14328 36139 14331
rect 36909 14331 36967 14337
rect 36909 14328 36921 14331
rect 36127 14300 36921 14328
rect 36127 14297 36139 14300
rect 36081 14291 36139 14297
rect 36909 14297 36921 14300
rect 36955 14297 36967 14331
rect 36909 14291 36967 14297
rect 28902 14260 28908 14272
rect 27948 14232 28396 14260
rect 28863 14232 28908 14260
rect 27948 14220 27954 14232
rect 28902 14220 28908 14232
rect 28960 14220 28966 14272
rect 33870 14220 33876 14272
rect 33928 14220 33934 14272
rect 33962 14220 33968 14272
rect 34020 14260 34026 14272
rect 34422 14260 34428 14272
rect 34020 14232 34428 14260
rect 34020 14220 34026 14232
rect 34422 14220 34428 14232
rect 34480 14260 34486 14272
rect 36096 14260 36124 14291
rect 36998 14288 37004 14340
rect 37056 14328 37062 14340
rect 37752 14328 37780 14359
rect 38378 14356 38384 14408
rect 38436 14396 38442 14408
rect 38565 14399 38623 14405
rect 38565 14396 38577 14399
rect 38436 14368 38577 14396
rect 38436 14356 38442 14368
rect 38565 14365 38577 14368
rect 38611 14365 38623 14399
rect 38565 14359 38623 14365
rect 38654 14356 38660 14408
rect 38712 14396 38718 14408
rect 38841 14399 38899 14405
rect 38841 14396 38853 14399
rect 38712 14368 38853 14396
rect 38712 14356 38718 14368
rect 38841 14365 38853 14368
rect 38887 14365 38899 14399
rect 38841 14359 38899 14365
rect 39025 14399 39083 14405
rect 39025 14365 39037 14399
rect 39071 14365 39083 14399
rect 39025 14359 39083 14365
rect 37056 14300 37780 14328
rect 37056 14288 37062 14300
rect 38470 14288 38476 14340
rect 38528 14328 38534 14340
rect 39040 14328 39068 14359
rect 39942 14356 39948 14408
rect 40000 14396 40006 14408
rect 40313 14399 40371 14405
rect 40313 14396 40325 14399
rect 40000 14368 40325 14396
rect 40000 14356 40006 14368
rect 40313 14365 40325 14368
rect 40359 14365 40371 14399
rect 40313 14359 40371 14365
rect 41601 14399 41659 14405
rect 41601 14365 41613 14399
rect 41647 14396 41659 14399
rect 41690 14396 41696 14408
rect 41647 14368 41696 14396
rect 41647 14365 41659 14368
rect 41601 14359 41659 14365
rect 41690 14356 41696 14368
rect 41748 14356 41754 14408
rect 41892 14405 41920 14572
rect 43070 14560 43076 14572
rect 43128 14600 43134 14612
rect 43717 14603 43775 14609
rect 43717 14600 43729 14603
rect 43128 14572 43729 14600
rect 43128 14560 43134 14572
rect 43717 14569 43729 14572
rect 43763 14569 43775 14603
rect 44453 14603 44511 14609
rect 44453 14600 44465 14603
rect 43717 14563 43775 14569
rect 43824 14572 44465 14600
rect 42613 14535 42671 14541
rect 42613 14501 42625 14535
rect 42659 14532 42671 14535
rect 43254 14532 43260 14544
rect 42659 14504 43260 14532
rect 42659 14501 42671 14504
rect 42613 14495 42671 14501
rect 43254 14492 43260 14504
rect 43312 14492 43318 14544
rect 42705 14467 42763 14473
rect 42705 14433 42717 14467
rect 42751 14464 42763 14467
rect 43824 14464 43852 14572
rect 44453 14569 44465 14572
rect 44499 14600 44511 14603
rect 44910 14600 44916 14612
rect 44499 14572 44916 14600
rect 44499 14569 44511 14572
rect 44453 14563 44511 14569
rect 44910 14560 44916 14572
rect 44968 14560 44974 14612
rect 45554 14600 45560 14612
rect 45020 14572 45560 14600
rect 44174 14492 44180 14544
rect 44232 14532 44238 14544
rect 45020 14532 45048 14572
rect 45554 14560 45560 14572
rect 45612 14560 45618 14612
rect 45646 14560 45652 14612
rect 45704 14600 45710 14612
rect 45704 14572 45749 14600
rect 45704 14560 45710 14572
rect 46014 14560 46020 14612
rect 46072 14600 46078 14612
rect 46845 14603 46903 14609
rect 46072 14560 46079 14600
rect 46845 14569 46857 14603
rect 46891 14600 46903 14603
rect 46934 14600 46940 14612
rect 46891 14572 46940 14600
rect 46891 14569 46903 14572
rect 46845 14563 46903 14569
rect 46934 14560 46940 14572
rect 46992 14560 46998 14612
rect 48038 14600 48044 14612
rect 47999 14572 48044 14600
rect 48038 14560 48044 14572
rect 48096 14560 48102 14612
rect 48148 14572 48820 14600
rect 44232 14504 45048 14532
rect 44232 14492 44238 14504
rect 45830 14492 45836 14544
rect 45888 14492 45894 14544
rect 42751 14436 43852 14464
rect 45848 14464 45876 14492
rect 45848 14436 45922 14464
rect 42751 14433 42763 14436
rect 42705 14427 42763 14433
rect 41877 14399 41935 14405
rect 41877 14365 41889 14399
rect 41923 14365 41935 14399
rect 42429 14399 42487 14405
rect 42429 14396 42441 14399
rect 41877 14359 41935 14365
rect 41984 14368 42441 14396
rect 38528 14300 39068 14328
rect 38528 14288 38534 14300
rect 41984 14272 42012 14368
rect 42429 14365 42441 14368
rect 42475 14365 42487 14399
rect 42429 14359 42487 14365
rect 42518 14356 42524 14408
rect 42576 14396 42582 14408
rect 42797 14399 42855 14405
rect 42576 14368 42621 14396
rect 42576 14356 42582 14368
rect 42797 14365 42809 14399
rect 42843 14396 42855 14399
rect 43898 14396 43904 14408
rect 42843 14368 43904 14396
rect 42843 14365 42855 14368
rect 42797 14359 42855 14365
rect 43898 14356 43904 14368
rect 43956 14356 43962 14408
rect 45646 14356 45652 14408
rect 45704 14396 45710 14408
rect 45894 14405 45922 14436
rect 46051 14405 46079 14560
rect 46290 14492 46296 14544
rect 46348 14532 46354 14544
rect 48148 14532 48176 14572
rect 46348 14504 48176 14532
rect 46348 14492 46354 14504
rect 48682 14492 48688 14544
rect 48740 14492 48746 14544
rect 48792 14532 48820 14572
rect 48866 14560 48872 14612
rect 48924 14600 48930 14612
rect 48961 14603 49019 14609
rect 48961 14600 48973 14603
rect 48924 14572 48973 14600
rect 48924 14560 48930 14572
rect 48961 14569 48973 14572
rect 49007 14569 49019 14603
rect 50614 14600 50620 14612
rect 48961 14563 49019 14569
rect 49620 14572 50620 14600
rect 49620 14532 49648 14572
rect 50614 14560 50620 14572
rect 50672 14560 50678 14612
rect 51166 14600 51172 14612
rect 51127 14572 51172 14600
rect 51166 14560 51172 14572
rect 51224 14560 51230 14612
rect 51902 14560 51908 14612
rect 51960 14600 51966 14612
rect 52178 14600 52184 14612
rect 51960 14572 52184 14600
rect 51960 14560 51966 14572
rect 52178 14560 52184 14572
rect 52236 14560 52242 14612
rect 52546 14600 52552 14612
rect 52507 14572 52552 14600
rect 52546 14560 52552 14572
rect 52604 14560 52610 14612
rect 52914 14560 52920 14612
rect 52972 14600 52978 14612
rect 53009 14603 53067 14609
rect 53009 14600 53021 14603
rect 52972 14572 53021 14600
rect 52972 14560 52978 14572
rect 53009 14569 53021 14572
rect 53055 14569 53067 14603
rect 54386 14600 54392 14612
rect 54347 14572 54392 14600
rect 53009 14563 53067 14569
rect 54386 14560 54392 14572
rect 54444 14560 54450 14612
rect 55122 14560 55128 14612
rect 55180 14600 55186 14612
rect 56226 14600 56232 14612
rect 55180 14572 56232 14600
rect 55180 14560 55186 14572
rect 56226 14560 56232 14572
rect 56284 14560 56290 14612
rect 57333 14603 57391 14609
rect 57333 14569 57345 14603
rect 57379 14600 57391 14603
rect 57606 14600 57612 14612
rect 57379 14572 57612 14600
rect 57379 14569 57391 14572
rect 57333 14563 57391 14569
rect 57606 14560 57612 14572
rect 57664 14560 57670 14612
rect 49786 14532 49792 14544
rect 48792 14504 49648 14532
rect 49747 14504 49792 14532
rect 49786 14492 49792 14504
rect 49844 14532 49850 14544
rect 49844 14504 50108 14532
rect 49844 14492 49850 14504
rect 46658 14424 46664 14476
rect 46716 14464 46722 14476
rect 48700 14464 48728 14492
rect 49970 14464 49976 14476
rect 46716 14436 47992 14464
rect 48700 14436 49976 14464
rect 46716 14424 46722 14436
rect 45879 14399 45937 14405
rect 45879 14396 45891 14399
rect 45704 14368 45891 14396
rect 45704 14356 45710 14368
rect 45879 14365 45891 14368
rect 45925 14365 45937 14399
rect 45879 14359 45937 14365
rect 46030 14399 46088 14405
rect 46293 14399 46351 14405
rect 46030 14365 46042 14399
rect 46076 14365 46088 14399
rect 46030 14359 46088 14365
rect 46130 14393 46188 14399
rect 46130 14359 46142 14393
rect 46176 14359 46188 14393
rect 46293 14365 46305 14399
rect 46339 14365 46351 14399
rect 47026 14396 47032 14408
rect 46987 14368 47032 14396
rect 46293 14359 46351 14365
rect 46130 14353 46188 14359
rect 43533 14331 43591 14337
rect 43533 14297 43545 14331
rect 43579 14328 43591 14331
rect 44174 14328 44180 14340
rect 43579 14300 44180 14328
rect 43579 14297 43591 14300
rect 43533 14291 43591 14297
rect 44174 14288 44180 14300
rect 44232 14328 44238 14340
rect 45370 14328 45376 14340
rect 44232 14300 45376 14328
rect 44232 14288 44238 14300
rect 45370 14288 45376 14300
rect 45428 14288 45434 14340
rect 34480 14232 36124 14260
rect 34480 14220 34486 14232
rect 36170 14220 36176 14272
rect 36228 14260 36234 14272
rect 36722 14269 36728 14272
rect 36709 14263 36728 14269
rect 36709 14260 36721 14263
rect 36228 14232 36721 14260
rect 36228 14220 36234 14232
rect 36709 14229 36721 14232
rect 36780 14260 36786 14272
rect 38194 14260 38200 14272
rect 36780 14232 38200 14260
rect 36709 14223 36728 14229
rect 36722 14220 36728 14223
rect 36780 14220 36786 14232
rect 38194 14220 38200 14232
rect 38252 14220 38258 14272
rect 41785 14263 41843 14269
rect 41785 14229 41797 14263
rect 41831 14260 41843 14263
rect 41966 14260 41972 14272
rect 41831 14232 41972 14260
rect 41831 14229 41843 14232
rect 41785 14223 41843 14229
rect 41966 14220 41972 14232
rect 42024 14220 42030 14272
rect 43438 14220 43444 14272
rect 43496 14260 43502 14272
rect 43733 14263 43791 14269
rect 43733 14260 43745 14263
rect 43496 14232 43745 14260
rect 43496 14220 43502 14232
rect 43733 14229 43745 14232
rect 43779 14229 43791 14263
rect 43733 14223 43791 14229
rect 43901 14263 43959 14269
rect 43901 14229 43913 14263
rect 43947 14260 43959 14263
rect 45554 14260 45560 14272
rect 43947 14232 45560 14260
rect 43947 14229 43959 14232
rect 43901 14223 43959 14229
rect 45554 14220 45560 14232
rect 45612 14220 45618 14272
rect 45738 14220 45744 14272
rect 45796 14260 45802 14272
rect 46144 14260 46172 14353
rect 46308 14272 46336 14359
rect 47026 14356 47032 14368
rect 47084 14356 47090 14408
rect 47118 14356 47124 14408
rect 47176 14396 47182 14408
rect 47394 14396 47400 14408
rect 47176 14368 47221 14396
rect 47355 14368 47400 14396
rect 47176 14356 47182 14368
rect 47394 14356 47400 14368
rect 47452 14356 47458 14408
rect 47489 14399 47547 14405
rect 47489 14365 47501 14399
rect 47535 14396 47547 14399
rect 47964 14396 47992 14436
rect 48225 14399 48283 14405
rect 48225 14396 48237 14399
rect 47535 14368 47900 14396
rect 47964 14368 48237 14396
rect 47535 14365 47547 14368
rect 47489 14359 47547 14365
rect 46934 14288 46940 14340
rect 46992 14328 46998 14340
rect 47213 14331 47271 14337
rect 47213 14328 47225 14331
rect 46992 14300 47225 14328
rect 46992 14288 46998 14300
rect 47213 14297 47225 14300
rect 47259 14328 47271 14331
rect 47762 14328 47768 14340
rect 47259 14300 47768 14328
rect 47259 14297 47271 14300
rect 47213 14291 47271 14297
rect 47762 14288 47768 14300
rect 47820 14288 47826 14340
rect 47872 14328 47900 14368
rect 48225 14365 48237 14368
rect 48271 14365 48283 14399
rect 48225 14359 48283 14365
rect 48406 14356 48412 14408
rect 48464 14356 48470 14408
rect 48501 14399 48559 14405
rect 48501 14365 48513 14399
rect 48547 14396 48559 14399
rect 48682 14396 48688 14408
rect 48547 14368 48688 14396
rect 48547 14365 48559 14368
rect 48501 14359 48559 14365
rect 48682 14356 48688 14368
rect 48740 14396 48746 14408
rect 49050 14396 49056 14408
rect 48740 14368 49056 14396
rect 48740 14356 48746 14368
rect 49050 14356 49056 14368
rect 49108 14356 49114 14408
rect 49160 14405 49188 14436
rect 49970 14424 49976 14436
rect 50028 14424 50034 14476
rect 49145 14399 49203 14405
rect 49145 14365 49157 14399
rect 49191 14365 49203 14399
rect 49145 14359 49203 14365
rect 49237 14399 49295 14405
rect 49237 14365 49249 14399
rect 49283 14396 49295 14399
rect 49326 14396 49332 14408
rect 49283 14368 49332 14396
rect 49283 14365 49295 14368
rect 49237 14359 49295 14365
rect 49326 14356 49332 14368
rect 49384 14356 49390 14408
rect 50080 14396 50108 14504
rect 50154 14492 50160 14544
rect 50212 14532 50218 14544
rect 50985 14535 51043 14541
rect 50985 14532 50997 14535
rect 50212 14504 50997 14532
rect 50212 14492 50218 14504
rect 50985 14501 50997 14504
rect 51031 14501 51043 14535
rect 50985 14495 51043 14501
rect 51077 14535 51135 14541
rect 51077 14501 51089 14535
rect 51123 14532 51135 14535
rect 53098 14532 53104 14544
rect 51123 14504 53104 14532
rect 51123 14501 51135 14504
rect 51077 14495 51135 14501
rect 53098 14492 53104 14504
rect 53156 14492 53162 14544
rect 50801 14467 50859 14473
rect 50801 14433 50813 14467
rect 50847 14464 50859 14467
rect 52181 14467 52239 14473
rect 52181 14464 52193 14467
rect 50847 14436 52193 14464
rect 50847 14433 50859 14436
rect 50801 14427 50859 14433
rect 52181 14433 52193 14436
rect 52227 14433 52239 14467
rect 52181 14427 52239 14433
rect 52638 14424 52644 14476
rect 52696 14464 52702 14476
rect 55585 14467 55643 14473
rect 55585 14464 55597 14467
rect 52696 14436 55597 14464
rect 52696 14424 52702 14436
rect 51166 14396 51172 14408
rect 50080 14368 51172 14396
rect 51166 14356 51172 14368
rect 51224 14396 51230 14408
rect 51261 14399 51319 14405
rect 51261 14396 51273 14399
rect 51224 14368 51273 14396
rect 51224 14356 51230 14368
rect 51261 14365 51273 14368
rect 51307 14365 51319 14399
rect 51902 14396 51908 14408
rect 51863 14368 51908 14396
rect 51261 14359 51319 14365
rect 51902 14356 51908 14368
rect 51960 14356 51966 14408
rect 52086 14396 52092 14408
rect 52047 14368 52092 14396
rect 52086 14356 52092 14368
rect 52144 14356 52150 14408
rect 52270 14396 52276 14408
rect 52231 14368 52276 14396
rect 52270 14356 52276 14368
rect 52328 14356 52334 14408
rect 52365 14399 52423 14405
rect 52365 14365 52377 14399
rect 52411 14396 52423 14399
rect 52454 14396 52460 14408
rect 52411 14368 52460 14396
rect 52411 14365 52423 14368
rect 52365 14359 52423 14365
rect 52454 14356 52460 14368
rect 52512 14396 52518 14408
rect 52730 14396 52736 14408
rect 52512 14368 52736 14396
rect 52512 14356 52518 14368
rect 52730 14356 52736 14368
rect 52788 14356 52794 14408
rect 53193 14399 53251 14405
rect 53193 14365 53205 14399
rect 53239 14365 53251 14399
rect 53193 14359 53251 14365
rect 48314 14328 48320 14340
rect 47872 14300 48320 14328
rect 46290 14260 46296 14272
rect 45796 14232 46172 14260
rect 46203 14232 46296 14260
rect 45796 14220 45802 14232
rect 46290 14220 46296 14232
rect 46348 14260 46354 14272
rect 47872 14260 47900 14300
rect 48314 14288 48320 14300
rect 48372 14288 48378 14340
rect 48424 14328 48452 14356
rect 48961 14331 49019 14337
rect 48961 14328 48973 14331
rect 48424 14300 48973 14328
rect 48961 14297 48973 14300
rect 49007 14328 49019 14331
rect 49007 14300 49740 14328
rect 49007 14297 49019 14300
rect 48961 14291 49019 14297
rect 46348 14232 47900 14260
rect 48409 14263 48467 14269
rect 46348 14220 46354 14232
rect 48409 14229 48421 14263
rect 48455 14260 48467 14263
rect 49050 14260 49056 14272
rect 48455 14232 49056 14260
rect 48455 14229 48467 14232
rect 48409 14223 48467 14229
rect 49050 14220 49056 14232
rect 49108 14220 49114 14272
rect 49712 14260 49740 14300
rect 51534 14288 51540 14340
rect 51592 14328 51598 14340
rect 53208 14328 53236 14359
rect 53282 14356 53288 14408
rect 53340 14396 53346 14408
rect 53484 14405 53512 14436
rect 53469 14399 53527 14405
rect 53340 14368 53385 14396
rect 53340 14356 53346 14368
rect 53469 14365 53481 14399
rect 53515 14365 53527 14399
rect 53469 14359 53527 14365
rect 53561 14399 53619 14405
rect 53561 14365 53573 14399
rect 53607 14365 53619 14399
rect 53561 14359 53619 14365
rect 53576 14328 53604 14359
rect 53834 14356 53840 14408
rect 53892 14396 53898 14408
rect 54220 14405 54248 14436
rect 55585 14433 55597 14436
rect 55631 14433 55643 14467
rect 55585 14427 55643 14433
rect 54021 14399 54079 14405
rect 54021 14396 54033 14399
rect 53892 14368 54033 14396
rect 53892 14356 53898 14368
rect 54021 14365 54033 14368
rect 54067 14365 54079 14399
rect 54021 14359 54079 14365
rect 54205 14399 54263 14405
rect 54205 14365 54217 14399
rect 54251 14365 54263 14399
rect 54205 14359 54263 14365
rect 54570 14356 54576 14408
rect 54628 14396 54634 14408
rect 55493 14399 55551 14405
rect 55493 14396 55505 14399
rect 54628 14368 55505 14396
rect 54628 14356 54634 14368
rect 55493 14365 55505 14368
rect 55539 14365 55551 14399
rect 55493 14359 55551 14365
rect 55674 14356 55680 14408
rect 55732 14396 55738 14408
rect 57882 14396 57888 14408
rect 55732 14368 57888 14396
rect 55732 14356 55738 14368
rect 57882 14356 57888 14368
rect 57940 14356 57946 14408
rect 51592 14300 53236 14328
rect 53392 14300 53604 14328
rect 51592 14288 51598 14300
rect 50338 14260 50344 14272
rect 49712 14232 50344 14260
rect 50338 14220 50344 14232
rect 50396 14220 50402 14272
rect 51353 14263 51411 14269
rect 51353 14229 51365 14263
rect 51399 14260 51411 14263
rect 52270 14260 52276 14272
rect 51399 14232 52276 14260
rect 51399 14229 51411 14232
rect 51353 14223 51411 14229
rect 52270 14220 52276 14232
rect 52328 14220 52334 14272
rect 53098 14220 53104 14272
rect 53156 14260 53162 14272
rect 53392 14260 53420 14300
rect 53156 14232 53420 14260
rect 53156 14220 53162 14232
rect 54386 14220 54392 14272
rect 54444 14260 54450 14272
rect 54846 14260 54852 14272
rect 54444 14232 54852 14260
rect 54444 14220 54450 14232
rect 54846 14220 54852 14232
rect 54904 14220 54910 14272
rect 56686 14260 56692 14272
rect 56647 14232 56692 14260
rect 56686 14220 56692 14232
rect 56744 14220 56750 14272
rect 57790 14260 57796 14272
rect 57751 14232 57796 14260
rect 57790 14220 57796 14232
rect 57848 14260 57854 14272
rect 58066 14260 58072 14272
rect 57848 14232 58072 14260
rect 57848 14220 57854 14232
rect 58066 14220 58072 14232
rect 58124 14220 58130 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 28718 14056 28724 14068
rect 24964 14028 28258 14056
rect 28679 14028 28724 14056
rect 24964 13932 24992 14028
rect 26237 13991 26295 13997
rect 26237 13957 26249 13991
rect 26283 13988 26295 13991
rect 26418 13988 26424 14000
rect 26283 13960 26424 13988
rect 26283 13957 26295 13960
rect 26237 13951 26295 13957
rect 26418 13948 26424 13960
rect 26476 13988 26482 14000
rect 27890 13988 27896 14000
rect 26476 13960 27896 13988
rect 26476 13948 26482 13960
rect 27890 13948 27896 13960
rect 27948 13988 27954 14000
rect 27948 13960 28028 13988
rect 27948 13948 27954 13960
rect 24946 13920 24952 13932
rect 24859 13892 24952 13920
rect 24946 13880 24952 13892
rect 25004 13880 25010 13932
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13920 25651 13923
rect 25774 13920 25780 13932
rect 25639 13892 25780 13920
rect 25639 13889 25651 13892
rect 25593 13883 25651 13889
rect 24213 13855 24271 13861
rect 24213 13821 24225 13855
rect 24259 13852 24271 13855
rect 25424 13852 25452 13883
rect 25774 13880 25780 13892
rect 25832 13920 25838 13932
rect 26142 13920 26148 13932
rect 25832 13892 26148 13920
rect 25832 13880 25838 13892
rect 26142 13880 26148 13892
rect 26200 13920 26206 13932
rect 26329 13923 26387 13929
rect 26329 13920 26341 13923
rect 26200 13892 26341 13920
rect 26200 13880 26206 13892
rect 26329 13889 26341 13892
rect 26375 13889 26387 13923
rect 26329 13883 26387 13889
rect 26510 13880 26516 13932
rect 26568 13920 26574 13932
rect 26605 13923 26663 13929
rect 26605 13920 26617 13923
rect 26568 13892 26617 13920
rect 26568 13880 26574 13892
rect 26605 13889 26617 13892
rect 26651 13920 26663 13923
rect 26970 13920 26976 13932
rect 26651 13892 26976 13920
rect 26651 13889 26663 13892
rect 26605 13883 26663 13889
rect 26970 13880 26976 13892
rect 27028 13880 27034 13932
rect 28000 13929 28028 13960
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13889 27859 13923
rect 27801 13883 27859 13889
rect 27985 13923 28043 13929
rect 27985 13889 27997 13923
rect 28031 13889 28043 13923
rect 27985 13883 28043 13889
rect 28077 13923 28135 13929
rect 28077 13889 28089 13923
rect 28123 13889 28135 13923
rect 28230 13920 28258 14028
rect 28718 14016 28724 14028
rect 28776 14016 28782 14068
rect 29365 14059 29423 14065
rect 29365 14025 29377 14059
rect 29411 14056 29423 14059
rect 30006 14056 30012 14068
rect 29411 14028 30012 14056
rect 29411 14025 29423 14028
rect 29365 14019 29423 14025
rect 30006 14016 30012 14028
rect 30064 14016 30070 14068
rect 30374 14016 30380 14068
rect 30432 14056 30438 14068
rect 30843 14059 30901 14065
rect 30843 14056 30855 14059
rect 30432 14028 30855 14056
rect 30432 14016 30438 14028
rect 30843 14025 30855 14028
rect 30889 14025 30901 14059
rect 31294 14056 31300 14068
rect 30843 14019 30901 14025
rect 30944 14028 31300 14056
rect 29730 13988 29736 14000
rect 29656 13960 29736 13988
rect 28629 13923 28687 13929
rect 28629 13920 28641 13923
rect 28230 13892 28641 13920
rect 28077 13883 28135 13889
rect 28629 13889 28641 13892
rect 28675 13889 28687 13923
rect 28810 13920 28816 13932
rect 28771 13892 28816 13920
rect 28629 13883 28687 13889
rect 24259 13824 26188 13852
rect 24259 13821 24271 13824
rect 24213 13815 24271 13821
rect 24765 13787 24823 13793
rect 24765 13753 24777 13787
rect 24811 13784 24823 13787
rect 25958 13784 25964 13796
rect 24811 13756 25964 13784
rect 24811 13753 24823 13756
rect 24765 13747 24823 13753
rect 25958 13744 25964 13756
rect 26016 13744 26022 13796
rect 26160 13784 26188 13824
rect 26234 13812 26240 13864
rect 26292 13852 26298 13864
rect 27617 13855 27675 13861
rect 27617 13852 27629 13855
rect 26292 13824 27629 13852
rect 26292 13812 26298 13824
rect 27617 13821 27629 13824
rect 27663 13821 27675 13855
rect 27617 13815 27675 13821
rect 26878 13784 26884 13796
rect 26160 13756 26884 13784
rect 26878 13744 26884 13756
rect 26936 13744 26942 13796
rect 25685 13719 25743 13725
rect 25685 13685 25697 13719
rect 25731 13716 25743 13719
rect 26050 13716 26056 13728
rect 25731 13688 26056 13716
rect 25731 13685 25743 13688
rect 25685 13679 25743 13685
rect 26050 13676 26056 13688
rect 26108 13676 26114 13728
rect 27816 13716 27844 13883
rect 27893 13855 27951 13861
rect 27893 13821 27905 13855
rect 27939 13821 27951 13855
rect 28092 13852 28120 13883
rect 28810 13880 28816 13892
rect 28868 13880 28874 13932
rect 29362 13920 29368 13932
rect 29323 13892 29368 13920
rect 29362 13880 29368 13892
rect 29420 13880 29426 13932
rect 29546 13920 29552 13932
rect 29507 13892 29552 13920
rect 29546 13880 29552 13892
rect 29604 13880 29610 13932
rect 29656 13929 29684 13960
rect 29730 13948 29736 13960
rect 29788 13948 29794 14000
rect 30745 13991 30803 13997
rect 30745 13957 30757 13991
rect 30791 13988 30803 13991
rect 30944 13988 30972 14028
rect 31294 14016 31300 14028
rect 31352 14016 31358 14068
rect 32309 14059 32367 14065
rect 32309 14025 32321 14059
rect 32355 14056 32367 14059
rect 32490 14056 32496 14068
rect 32355 14028 32496 14056
rect 32355 14025 32367 14028
rect 32309 14019 32367 14025
rect 32490 14016 32496 14028
rect 32548 14016 32554 14068
rect 33594 14016 33600 14068
rect 33652 14016 33658 14068
rect 33686 14016 33692 14068
rect 33744 14056 33750 14068
rect 34517 14059 34575 14065
rect 34517 14056 34529 14059
rect 33744 14028 34529 14056
rect 33744 14016 33750 14028
rect 34517 14025 34529 14028
rect 34563 14025 34575 14059
rect 34517 14019 34575 14025
rect 35621 14059 35679 14065
rect 35621 14025 35633 14059
rect 35667 14056 35679 14059
rect 35710 14056 35716 14068
rect 35667 14028 35716 14056
rect 35667 14025 35679 14028
rect 35621 14019 35679 14025
rect 35710 14016 35716 14028
rect 35768 14016 35774 14068
rect 36998 14056 37004 14068
rect 35912 14028 37004 14056
rect 33612 13988 33640 14016
rect 34885 13991 34943 13997
rect 30791 13960 30972 13988
rect 32784 13960 34468 13988
rect 30791 13957 30803 13960
rect 30745 13951 30803 13957
rect 29641 13923 29699 13929
rect 29641 13889 29653 13923
rect 29687 13889 29699 13923
rect 29914 13920 29920 13932
rect 29875 13892 29920 13920
rect 29641 13883 29699 13889
rect 29914 13880 29920 13892
rect 29972 13920 29978 13932
rect 30929 13923 30987 13929
rect 30929 13920 30941 13923
rect 29972 13892 30941 13920
rect 29972 13880 29978 13892
rect 30929 13889 30941 13892
rect 30975 13889 30987 13923
rect 30929 13883 30987 13889
rect 31018 13880 31024 13932
rect 31076 13920 31082 13932
rect 31076 13892 31121 13920
rect 31076 13880 31082 13892
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 32493 13923 32551 13929
rect 32493 13920 32505 13923
rect 31720 13892 32505 13920
rect 31720 13880 31726 13892
rect 32493 13889 32505 13892
rect 32539 13889 32551 13923
rect 32493 13883 32551 13889
rect 32582 13880 32588 13932
rect 32640 13920 32646 13932
rect 32784 13929 32812 13960
rect 32677 13923 32735 13929
rect 32677 13920 32689 13923
rect 32640 13892 32689 13920
rect 32640 13880 32646 13892
rect 32677 13889 32689 13892
rect 32723 13889 32735 13923
rect 32677 13883 32735 13889
rect 32769 13923 32827 13929
rect 32769 13889 32781 13923
rect 32815 13889 32827 13923
rect 32769 13883 32827 13889
rect 32950 13880 32956 13932
rect 33008 13920 33014 13932
rect 33229 13923 33287 13929
rect 33229 13920 33241 13923
rect 33008 13892 33241 13920
rect 33008 13880 33014 13892
rect 33229 13889 33241 13892
rect 33275 13889 33287 13923
rect 33410 13920 33416 13932
rect 33371 13892 33416 13920
rect 33229 13883 33287 13889
rect 33410 13880 33416 13892
rect 33468 13880 33474 13932
rect 33505 13923 33563 13929
rect 33505 13889 33517 13923
rect 33551 13889 33563 13923
rect 33505 13883 33563 13889
rect 33633 13923 33691 13929
rect 33633 13889 33645 13923
rect 33679 13920 33691 13923
rect 33870 13920 33876 13932
rect 33679 13892 33876 13920
rect 33679 13889 33691 13892
rect 33633 13883 33691 13889
rect 28718 13852 28724 13864
rect 28092 13824 28724 13852
rect 27893 13815 27951 13821
rect 27908 13784 27936 13815
rect 28718 13812 28724 13824
rect 28776 13812 28782 13864
rect 29825 13855 29883 13861
rect 29825 13821 29837 13855
rect 29871 13852 29883 13855
rect 31754 13852 31760 13864
rect 29871 13824 31760 13852
rect 29871 13821 29883 13824
rect 29825 13815 29883 13821
rect 31754 13812 31760 13824
rect 31812 13852 31818 13864
rect 32214 13852 32220 13864
rect 31812 13824 32220 13852
rect 31812 13812 31818 13824
rect 32214 13812 32220 13824
rect 32272 13812 32278 13864
rect 33318 13852 33324 13864
rect 33279 13824 33324 13852
rect 33318 13812 33324 13824
rect 33376 13812 33382 13864
rect 33520 13852 33548 13883
rect 33870 13880 33876 13892
rect 33928 13880 33934 13932
rect 34440 13929 34468 13960
rect 34885 13957 34897 13991
rect 34931 13988 34943 13991
rect 35912 13988 35940 14028
rect 36998 14016 37004 14028
rect 37056 14016 37062 14068
rect 37274 14016 37280 14068
rect 37332 14056 37338 14068
rect 37461 14059 37519 14065
rect 37461 14056 37473 14059
rect 37332 14028 37473 14056
rect 37332 14016 37338 14028
rect 37461 14025 37473 14028
rect 37507 14025 37519 14059
rect 37461 14019 37519 14025
rect 38565 14059 38623 14065
rect 38565 14025 38577 14059
rect 38611 14056 38623 14059
rect 38654 14056 38660 14068
rect 38611 14028 38660 14056
rect 38611 14025 38623 14028
rect 38565 14019 38623 14025
rect 38654 14016 38660 14028
rect 38712 14016 38718 14068
rect 38749 14059 38807 14065
rect 38749 14025 38761 14059
rect 38795 14056 38807 14059
rect 38838 14056 38844 14068
rect 38795 14028 38844 14056
rect 38795 14025 38807 14028
rect 38749 14019 38807 14025
rect 38838 14016 38844 14028
rect 38896 14016 38902 14068
rect 41598 14056 41604 14068
rect 41559 14028 41604 14056
rect 41598 14016 41604 14028
rect 41656 14016 41662 14068
rect 43530 14016 43536 14068
rect 43588 14056 43594 14068
rect 43625 14059 43683 14065
rect 43625 14056 43637 14059
rect 43588 14028 43637 14056
rect 43588 14016 43594 14028
rect 43625 14025 43637 14028
rect 43671 14025 43683 14059
rect 43625 14019 43683 14025
rect 45465 14059 45523 14065
rect 45465 14025 45477 14059
rect 45511 14056 45523 14059
rect 45511 14028 45784 14056
rect 45511 14025 45523 14028
rect 45465 14019 45523 14025
rect 34931 13960 35940 13988
rect 35989 13991 36047 13997
rect 34931 13957 34943 13960
rect 34885 13951 34943 13957
rect 35989 13957 36001 13991
rect 36035 13988 36047 13991
rect 37366 13988 37372 14000
rect 36035 13960 37372 13988
rect 36035 13957 36047 13960
rect 35989 13951 36047 13957
rect 37366 13948 37372 13960
rect 37424 13948 37430 14000
rect 38470 13948 38476 14000
rect 38528 13988 38534 14000
rect 38528 13960 40080 13988
rect 38528 13948 38534 13960
rect 34425 13923 34483 13929
rect 34425 13889 34437 13923
rect 34471 13920 34483 13923
rect 34514 13920 34520 13932
rect 34471 13892 34520 13920
rect 34471 13889 34483 13892
rect 34425 13883 34483 13889
rect 34514 13880 34520 13892
rect 34572 13880 34578 13932
rect 34698 13880 34704 13932
rect 34756 13920 34762 13932
rect 35434 13920 35440 13932
rect 34756 13892 35440 13920
rect 34756 13880 34762 13892
rect 35434 13880 35440 13892
rect 35492 13880 35498 13932
rect 35802 13920 35808 13932
rect 35763 13892 35808 13920
rect 35802 13880 35808 13892
rect 35860 13880 35866 13932
rect 35897 13923 35955 13929
rect 35897 13889 35909 13923
rect 35943 13889 35955 13923
rect 35897 13883 35955 13889
rect 36173 13923 36231 13929
rect 36173 13889 36185 13923
rect 36219 13889 36231 13923
rect 36173 13883 36231 13889
rect 35912 13852 35940 13883
rect 36078 13852 36084 13864
rect 33520 13824 36084 13852
rect 36078 13812 36084 13824
rect 36136 13812 36142 13864
rect 36188 13852 36216 13883
rect 36262 13880 36268 13932
rect 36320 13920 36326 13932
rect 36725 13923 36783 13929
rect 36725 13920 36737 13923
rect 36320 13892 36737 13920
rect 36320 13880 36326 13892
rect 36725 13889 36737 13892
rect 36771 13889 36783 13923
rect 36906 13920 36912 13932
rect 36867 13892 36912 13920
rect 36725 13883 36783 13889
rect 36354 13852 36360 13864
rect 36188 13824 36360 13852
rect 36354 13812 36360 13824
rect 36412 13812 36418 13864
rect 28902 13784 28908 13796
rect 27908 13756 28908 13784
rect 28902 13744 28908 13756
rect 28960 13784 28966 13796
rect 33502 13784 33508 13796
rect 28960 13756 29776 13784
rect 28960 13744 28966 13756
rect 29454 13716 29460 13728
rect 27816 13688 29460 13716
rect 29454 13676 29460 13688
rect 29512 13676 29518 13728
rect 29748 13716 29776 13756
rect 30852 13756 33508 13784
rect 30852 13716 30880 13756
rect 33502 13744 33508 13756
rect 33560 13744 33566 13796
rect 36740 13784 36768 13883
rect 36906 13880 36912 13892
rect 36964 13920 36970 13932
rect 37645 13923 37703 13929
rect 37645 13920 37657 13923
rect 36964 13892 37657 13920
rect 36964 13880 36970 13892
rect 37645 13889 37657 13892
rect 37691 13889 37703 13923
rect 37645 13883 37703 13889
rect 38746 13923 38804 13929
rect 38746 13889 38758 13923
rect 38792 13889 38804 13923
rect 39206 13920 39212 13932
rect 39167 13892 39212 13920
rect 38746 13883 38804 13889
rect 36817 13855 36875 13861
rect 36817 13821 36829 13855
rect 36863 13852 36875 13855
rect 37182 13852 37188 13864
rect 36863 13824 37188 13852
rect 36863 13821 36875 13824
rect 36817 13815 36875 13821
rect 37182 13812 37188 13824
rect 37240 13812 37246 13864
rect 37829 13855 37887 13861
rect 37829 13821 37841 13855
rect 37875 13821 37887 13855
rect 38761 13852 38789 13883
rect 39206 13880 39212 13892
rect 39264 13880 39270 13932
rect 39850 13920 39856 13932
rect 39811 13892 39856 13920
rect 39850 13880 39856 13892
rect 39908 13880 39914 13932
rect 40052 13929 40080 13960
rect 42978 13948 42984 14000
rect 43036 13988 43042 14000
rect 43441 13991 43499 13997
rect 43441 13988 43453 13991
rect 43036 13960 43453 13988
rect 43036 13948 43042 13960
rect 43441 13957 43453 13960
rect 43487 13957 43499 13991
rect 43441 13951 43499 13957
rect 43548 13960 45692 13988
rect 40037 13923 40095 13929
rect 40037 13889 40049 13923
rect 40083 13889 40095 13923
rect 40494 13920 40500 13932
rect 40455 13892 40500 13920
rect 40037 13883 40095 13889
rect 40494 13880 40500 13892
rect 40552 13880 40558 13932
rect 41417 13923 41475 13929
rect 41417 13889 41429 13923
rect 41463 13889 41475 13923
rect 41417 13883 41475 13889
rect 42705 13923 42763 13929
rect 42705 13889 42717 13923
rect 42751 13920 42763 13923
rect 43257 13923 43315 13929
rect 43257 13920 43269 13923
rect 42751 13892 43269 13920
rect 42751 13889 42763 13892
rect 42705 13883 42763 13889
rect 43257 13889 43269 13892
rect 43303 13920 43315 13923
rect 43346 13920 43352 13932
rect 43303 13892 43352 13920
rect 43303 13889 43315 13892
rect 43257 13883 43315 13889
rect 39114 13852 39120 13864
rect 38761 13824 39120 13852
rect 37829 13815 37887 13821
rect 37844 13784 37872 13815
rect 39114 13812 39120 13824
rect 39172 13852 39178 13864
rect 39868 13852 39896 13880
rect 39172 13824 39896 13852
rect 39945 13855 40003 13861
rect 39172 13812 39178 13824
rect 39945 13821 39957 13855
rect 39991 13852 40003 13855
rect 40402 13852 40408 13864
rect 39991 13824 40408 13852
rect 39991 13821 40003 13824
rect 39945 13815 40003 13821
rect 40402 13812 40408 13824
rect 40460 13812 40466 13864
rect 40957 13855 41015 13861
rect 40957 13821 40969 13855
rect 41003 13852 41015 13855
rect 41432 13852 41460 13883
rect 43346 13880 43352 13892
rect 43404 13880 43410 13932
rect 41003 13824 41460 13852
rect 41003 13821 41015 13824
rect 40957 13815 41015 13821
rect 41690 13812 41696 13864
rect 41748 13852 41754 13864
rect 42334 13852 42340 13864
rect 41748 13824 42340 13852
rect 41748 13812 41754 13824
rect 42334 13812 42340 13824
rect 42392 13852 42398 13864
rect 43548 13852 43576 13960
rect 44358 13880 44364 13932
rect 44416 13920 44422 13932
rect 44542 13920 44548 13932
rect 44416 13892 44548 13920
rect 44416 13880 44422 13892
rect 44542 13880 44548 13892
rect 44600 13880 44606 13932
rect 44729 13923 44787 13929
rect 44729 13889 44741 13923
rect 44775 13920 44787 13923
rect 45278 13920 45284 13932
rect 44775 13892 45284 13920
rect 44775 13889 44787 13892
rect 44729 13883 44787 13889
rect 45278 13880 45284 13892
rect 45336 13880 45342 13932
rect 45370 13880 45376 13932
rect 45428 13920 45434 13932
rect 45557 13923 45615 13929
rect 45428 13892 45473 13920
rect 45428 13880 45434 13892
rect 45557 13889 45569 13923
rect 45603 13889 45615 13923
rect 45557 13883 45615 13889
rect 42392 13824 43576 13852
rect 42392 13812 42398 13824
rect 44818 13812 44824 13864
rect 44876 13852 44882 13864
rect 45572 13852 45600 13883
rect 44876 13824 45600 13852
rect 45664 13852 45692 13960
rect 45756 13920 45784 14028
rect 45922 14016 45928 14068
rect 45980 14056 45986 14068
rect 46842 14056 46848 14068
rect 45980 14028 46848 14056
rect 45980 14016 45986 14028
rect 46842 14016 46848 14028
rect 46900 14056 46906 14068
rect 47026 14056 47032 14068
rect 46900 14028 47032 14056
rect 46900 14016 46906 14028
rect 47026 14016 47032 14028
rect 47084 14016 47090 14068
rect 47213 14059 47271 14065
rect 47213 14025 47225 14059
rect 47259 14056 47271 14059
rect 47394 14056 47400 14068
rect 47259 14028 47400 14056
rect 47259 14025 47271 14028
rect 47213 14019 47271 14025
rect 47394 14016 47400 14028
rect 47452 14016 47458 14068
rect 47854 14016 47860 14068
rect 47912 14056 47918 14068
rect 50617 14059 50675 14065
rect 47912 14028 50292 14056
rect 47912 14016 47918 14028
rect 50154 13988 50160 14000
rect 46400 13960 50160 13988
rect 45830 13920 45836 13932
rect 45743 13892 45836 13920
rect 45830 13880 45836 13892
rect 45888 13920 45894 13932
rect 46198 13920 46204 13932
rect 45888 13892 46204 13920
rect 45888 13880 45894 13892
rect 46198 13880 46204 13892
rect 46256 13880 46262 13932
rect 46400 13852 46428 13960
rect 50154 13948 50160 13960
rect 50212 13948 50218 14000
rect 50264 13988 50292 14028
rect 50617 14025 50629 14059
rect 50663 14025 50675 14059
rect 50617 14019 50675 14025
rect 51169 14059 51227 14065
rect 51169 14025 51181 14059
rect 51215 14056 51227 14059
rect 52086 14056 52092 14068
rect 51215 14028 52092 14056
rect 51215 14025 51227 14028
rect 51169 14019 51227 14025
rect 50632 13988 50660 14019
rect 52086 14016 52092 14028
rect 52144 14016 52150 14068
rect 52273 14059 52331 14065
rect 52273 14025 52285 14059
rect 52319 14056 52331 14059
rect 52362 14056 52368 14068
rect 52319 14028 52368 14056
rect 52319 14025 52331 14028
rect 52273 14019 52331 14025
rect 52362 14016 52368 14028
rect 52420 14016 52426 14068
rect 53374 14016 53380 14068
rect 53432 14056 53438 14068
rect 53561 14059 53619 14065
rect 53561 14056 53573 14059
rect 53432 14028 53573 14056
rect 53432 14016 53438 14028
rect 53561 14025 53573 14028
rect 53607 14025 53619 14059
rect 53561 14019 53619 14025
rect 54481 14059 54539 14065
rect 54481 14025 54493 14059
rect 54527 14056 54539 14059
rect 54662 14056 54668 14068
rect 54527 14028 54668 14056
rect 54527 14025 54539 14028
rect 54481 14019 54539 14025
rect 54662 14016 54668 14028
rect 54720 14016 54726 14068
rect 55122 14056 55128 14068
rect 55083 14028 55128 14056
rect 55122 14016 55128 14028
rect 55180 14016 55186 14068
rect 55214 14016 55220 14068
rect 55272 14056 55278 14068
rect 56226 14056 56232 14068
rect 55272 14028 56232 14056
rect 55272 14016 55278 14028
rect 51534 13988 51540 14000
rect 50264 13960 50384 13988
rect 50632 13960 51540 13988
rect 46477 13923 46535 13929
rect 46477 13889 46489 13923
rect 46523 13889 46535 13923
rect 46658 13920 46664 13932
rect 46619 13892 46664 13920
rect 46477 13883 46535 13889
rect 45664 13824 46428 13852
rect 44876 13812 44882 13824
rect 38470 13784 38476 13796
rect 36740 13756 38476 13784
rect 38470 13744 38476 13756
rect 38528 13744 38534 13796
rect 43530 13744 43536 13796
rect 43588 13784 43594 13796
rect 44836 13784 44864 13812
rect 43588 13756 44864 13784
rect 43588 13744 43594 13756
rect 29748 13688 30880 13716
rect 31110 13676 31116 13728
rect 31168 13716 31174 13728
rect 32122 13716 32128 13728
rect 31168 13688 32128 13716
rect 31168 13676 31174 13688
rect 32122 13676 32128 13688
rect 32180 13716 32186 13728
rect 37918 13716 37924 13728
rect 32180 13688 37924 13716
rect 32180 13676 32186 13688
rect 37918 13676 37924 13688
rect 37976 13676 37982 13728
rect 39117 13719 39175 13725
rect 39117 13685 39129 13719
rect 39163 13716 39175 13719
rect 39206 13716 39212 13728
rect 39163 13688 39212 13716
rect 39163 13685 39175 13688
rect 39117 13679 39175 13685
rect 39206 13676 39212 13688
rect 39264 13676 39270 13728
rect 40218 13676 40224 13728
rect 40276 13716 40282 13728
rect 40589 13719 40647 13725
rect 40589 13716 40601 13719
rect 40276 13688 40601 13716
rect 40276 13676 40282 13688
rect 40589 13685 40601 13688
rect 40635 13685 40647 13719
rect 44634 13716 44640 13728
rect 44595 13688 44640 13716
rect 40589 13679 40647 13685
rect 44634 13676 44640 13688
rect 44692 13676 44698 13728
rect 46492 13716 46520 13883
rect 46658 13880 46664 13892
rect 46716 13880 46722 13932
rect 46842 13920 46848 13932
rect 46803 13892 46848 13920
rect 46842 13880 46848 13892
rect 46900 13880 46906 13932
rect 47029 13923 47087 13929
rect 47029 13889 47041 13923
rect 47075 13920 47087 13923
rect 47394 13920 47400 13932
rect 47075 13892 47400 13920
rect 47075 13889 47087 13892
rect 47029 13883 47087 13889
rect 47394 13880 47400 13892
rect 47452 13880 47458 13932
rect 48498 13880 48504 13932
rect 48556 13920 48562 13932
rect 48777 13923 48835 13929
rect 48777 13920 48789 13923
rect 48556 13892 48789 13920
rect 48556 13880 48562 13892
rect 48777 13889 48789 13892
rect 48823 13889 48835 13923
rect 48777 13883 48835 13889
rect 48961 13923 49019 13929
rect 48961 13889 48973 13923
rect 49007 13889 49019 13923
rect 48961 13883 49019 13889
rect 46750 13852 46756 13864
rect 46711 13824 46756 13852
rect 46750 13812 46756 13824
rect 46808 13812 46814 13864
rect 47762 13852 47768 13864
rect 47723 13824 47768 13852
rect 47762 13812 47768 13824
rect 47820 13812 47826 13864
rect 48976 13728 49004 13883
rect 49145 13855 49203 13861
rect 49145 13821 49157 13855
rect 49191 13852 49203 13855
rect 49418 13852 49424 13864
rect 49191 13824 49424 13852
rect 49191 13821 49203 13824
rect 49145 13815 49203 13821
rect 49418 13812 49424 13824
rect 49476 13852 49482 13864
rect 49970 13852 49976 13864
rect 49476 13824 49976 13852
rect 49476 13812 49482 13824
rect 49970 13812 49976 13824
rect 50028 13812 50034 13864
rect 50154 13852 50160 13864
rect 50115 13824 50160 13852
rect 50154 13812 50160 13824
rect 50212 13812 50218 13864
rect 50356 13861 50384 13960
rect 51534 13948 51540 13960
rect 51592 13948 51598 14000
rect 53193 13991 53251 13997
rect 53193 13957 53205 13991
rect 53239 13988 53251 13991
rect 54846 13988 54852 14000
rect 53239 13960 54852 13988
rect 53239 13957 53251 13960
rect 53193 13951 53251 13957
rect 54846 13948 54852 13960
rect 54904 13948 54910 14000
rect 55490 13948 55496 14000
rect 55548 13988 55554 14000
rect 55677 13991 55735 13997
rect 55677 13988 55689 13991
rect 55548 13960 55689 13988
rect 55548 13948 55554 13960
rect 55677 13957 55689 13960
rect 55723 13957 55735 13991
rect 55677 13951 55735 13957
rect 50614 13880 50620 13932
rect 50672 13920 50678 13932
rect 51077 13923 51135 13929
rect 51077 13920 51089 13923
rect 50672 13892 51089 13920
rect 50672 13880 50678 13892
rect 51077 13889 51089 13892
rect 51123 13889 51135 13923
rect 51258 13920 51264 13932
rect 51219 13892 51264 13920
rect 51077 13883 51135 13889
rect 51258 13880 51264 13892
rect 51316 13880 51322 13932
rect 51626 13880 51632 13932
rect 51684 13920 51690 13932
rect 52181 13923 52239 13929
rect 52181 13920 52193 13923
rect 51684 13892 52193 13920
rect 51684 13880 51690 13892
rect 52181 13889 52193 13892
rect 52227 13889 52239 13923
rect 52181 13883 52239 13889
rect 52270 13880 52276 13932
rect 52328 13920 52334 13932
rect 52365 13923 52423 13929
rect 52365 13920 52377 13923
rect 52328 13892 52377 13920
rect 52328 13880 52334 13892
rect 52365 13889 52377 13892
rect 52411 13889 52423 13923
rect 52365 13883 52423 13889
rect 53101 13923 53159 13929
rect 53101 13889 53113 13923
rect 53147 13889 53159 13923
rect 53377 13923 53435 13929
rect 53377 13920 53389 13923
rect 53101 13883 53159 13889
rect 53300 13892 53389 13920
rect 50249 13855 50307 13861
rect 50249 13821 50261 13855
rect 50295 13821 50307 13855
rect 50249 13815 50307 13821
rect 50341 13855 50399 13861
rect 50341 13821 50353 13855
rect 50387 13821 50399 13855
rect 50341 13815 50399 13821
rect 49050 13744 49056 13796
rect 49108 13784 49114 13796
rect 50264 13784 50292 13815
rect 50430 13812 50436 13864
rect 50488 13852 50494 13864
rect 52822 13852 52828 13864
rect 50488 13824 50533 13852
rect 50632 13824 52828 13852
rect 50488 13812 50494 13824
rect 50632 13784 50660 13824
rect 52822 13812 52828 13824
rect 52880 13812 52886 13864
rect 49108 13756 50660 13784
rect 49108 13744 49114 13756
rect 51166 13744 51172 13796
rect 51224 13784 51230 13796
rect 52178 13784 52184 13796
rect 51224 13756 52184 13784
rect 51224 13744 51230 13756
rect 52178 13744 52184 13756
rect 52236 13784 52242 13796
rect 53116 13784 53144 13883
rect 53300 13864 53328 13892
rect 53377 13889 53389 13892
rect 53423 13889 53435 13923
rect 54202 13920 54208 13932
rect 54163 13892 54208 13920
rect 53377 13883 53435 13889
rect 54202 13880 54208 13892
rect 54260 13880 54266 13932
rect 54570 13920 54576 13932
rect 54531 13892 54576 13920
rect 54570 13880 54576 13892
rect 54628 13880 54634 13932
rect 55784 13929 55812 14028
rect 56226 14016 56232 14028
rect 56284 14056 56290 14068
rect 57606 14056 57612 14068
rect 56284 14028 57612 14056
rect 56284 14016 56290 14028
rect 57606 14016 57612 14028
rect 57664 14016 57670 14068
rect 58066 14056 58072 14068
rect 58027 14028 58072 14056
rect 58066 14016 58072 14028
rect 58124 14016 58130 14068
rect 57330 13988 57336 14000
rect 56704 13960 57336 13988
rect 55769 13923 55827 13929
rect 55769 13889 55781 13923
rect 55815 13889 55827 13923
rect 56042 13920 56048 13932
rect 56003 13892 56048 13920
rect 55769 13883 55827 13889
rect 56042 13880 56048 13892
rect 56100 13880 56106 13932
rect 56410 13880 56416 13932
rect 56468 13920 56474 13932
rect 56704 13929 56732 13960
rect 57330 13948 57336 13960
rect 57388 13948 57394 14000
rect 56689 13923 56747 13929
rect 56689 13920 56701 13923
rect 56468 13892 56701 13920
rect 56468 13880 56474 13892
rect 56689 13889 56701 13892
rect 56735 13889 56747 13923
rect 56689 13883 56747 13889
rect 56781 13923 56839 13929
rect 56781 13889 56793 13923
rect 56827 13889 56839 13923
rect 56781 13883 56839 13889
rect 53282 13812 53288 13864
rect 53340 13812 53346 13864
rect 53926 13812 53932 13864
rect 53984 13852 53990 13864
rect 54021 13855 54079 13861
rect 54021 13852 54033 13855
rect 53984 13824 54033 13852
rect 53984 13812 53990 13824
rect 54021 13821 54033 13824
rect 54067 13821 54079 13855
rect 54021 13815 54079 13821
rect 56502 13812 56508 13864
rect 56560 13852 56566 13864
rect 56796 13852 56824 13883
rect 56560 13824 56824 13852
rect 56560 13812 56566 13824
rect 53374 13784 53380 13796
rect 52236 13756 53380 13784
rect 52236 13744 52242 13756
rect 53374 13744 53380 13756
rect 53432 13784 53438 13796
rect 57790 13784 57796 13796
rect 53432 13756 57796 13784
rect 53432 13744 53438 13756
rect 57790 13744 57796 13756
rect 57848 13744 57854 13796
rect 48406 13716 48412 13728
rect 46492 13688 48412 13716
rect 48406 13676 48412 13688
rect 48464 13676 48470 13728
rect 48958 13676 48964 13728
rect 49016 13676 49022 13728
rect 49602 13676 49608 13728
rect 49660 13716 49666 13728
rect 52914 13716 52920 13728
rect 49660 13688 52920 13716
rect 49660 13676 49666 13688
rect 52914 13676 52920 13688
rect 52972 13676 52978 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 24946 13512 24952 13524
rect 24907 13484 24952 13512
rect 24946 13472 24952 13484
rect 25004 13472 25010 13524
rect 25682 13512 25688 13524
rect 25643 13484 25688 13512
rect 25682 13472 25688 13484
rect 25740 13472 25746 13524
rect 26053 13515 26111 13521
rect 26053 13481 26065 13515
rect 26099 13512 26111 13515
rect 26234 13512 26240 13524
rect 26099 13484 26240 13512
rect 26099 13481 26111 13484
rect 26053 13475 26111 13481
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 31294 13512 31300 13524
rect 28736 13484 31156 13512
rect 31255 13484 31300 13512
rect 26878 13404 26884 13456
rect 26936 13444 26942 13456
rect 27798 13444 27804 13456
rect 26936 13416 27804 13444
rect 26936 13404 26942 13416
rect 27798 13404 27804 13416
rect 27856 13404 27862 13456
rect 26050 13336 26056 13388
rect 26108 13376 26114 13388
rect 28736 13376 28764 13484
rect 31128 13444 31156 13484
rect 31294 13472 31300 13484
rect 31352 13472 31358 13524
rect 32122 13472 32128 13524
rect 32180 13512 32186 13524
rect 32309 13515 32367 13521
rect 32309 13512 32321 13515
rect 32180 13484 32321 13512
rect 32180 13472 32186 13484
rect 32309 13481 32321 13484
rect 32355 13481 32367 13515
rect 32309 13475 32367 13481
rect 33689 13515 33747 13521
rect 33689 13481 33701 13515
rect 33735 13512 33747 13515
rect 33870 13512 33876 13524
rect 33735 13484 33876 13512
rect 33735 13481 33747 13484
rect 33689 13475 33747 13481
rect 33870 13472 33876 13484
rect 33928 13472 33934 13524
rect 36081 13515 36139 13521
rect 36081 13481 36093 13515
rect 36127 13512 36139 13515
rect 36722 13512 36728 13524
rect 36127 13484 36728 13512
rect 36127 13481 36139 13484
rect 36081 13475 36139 13481
rect 36722 13472 36728 13484
rect 36780 13512 36786 13524
rect 37182 13512 37188 13524
rect 36780 13484 37188 13512
rect 36780 13472 36786 13484
rect 37182 13472 37188 13484
rect 37240 13472 37246 13524
rect 37366 13472 37372 13524
rect 37424 13512 37430 13524
rect 37461 13515 37519 13521
rect 37461 13512 37473 13515
rect 37424 13484 37473 13512
rect 37424 13472 37430 13484
rect 37461 13481 37473 13484
rect 37507 13481 37519 13515
rect 37461 13475 37519 13481
rect 38102 13472 38108 13524
rect 38160 13512 38166 13524
rect 39206 13512 39212 13524
rect 38160 13484 39212 13512
rect 38160 13472 38166 13484
rect 39206 13472 39212 13484
rect 39264 13472 39270 13524
rect 40037 13515 40095 13521
rect 40037 13481 40049 13515
rect 40083 13512 40095 13515
rect 40310 13512 40316 13524
rect 40083 13484 40316 13512
rect 40083 13481 40095 13484
rect 40037 13475 40095 13481
rect 40310 13472 40316 13484
rect 40368 13472 40374 13524
rect 43070 13512 43076 13524
rect 43031 13484 43076 13512
rect 43070 13472 43076 13484
rect 43128 13472 43134 13524
rect 44266 13512 44272 13524
rect 44227 13484 44272 13512
rect 44266 13472 44272 13484
rect 44324 13512 44330 13524
rect 46382 13512 46388 13524
rect 44324 13484 46244 13512
rect 46343 13484 46388 13512
rect 44324 13472 44330 13484
rect 31662 13444 31668 13456
rect 26108 13348 28764 13376
rect 28920 13416 30972 13444
rect 31128 13416 31668 13444
rect 26108 13336 26114 13348
rect 25866 13308 25872 13320
rect 25827 13280 25872 13308
rect 25866 13268 25872 13280
rect 25924 13268 25930 13320
rect 25958 13268 25964 13320
rect 26016 13308 26022 13320
rect 26145 13311 26203 13317
rect 26145 13308 26157 13311
rect 26016 13280 26157 13308
rect 26016 13268 26022 13280
rect 26145 13277 26157 13280
rect 26191 13277 26203 13311
rect 26878 13308 26884 13320
rect 26839 13280 26884 13308
rect 26145 13271 26203 13277
rect 26878 13268 26884 13280
rect 26936 13268 26942 13320
rect 27798 13308 27804 13320
rect 27759 13280 27804 13308
rect 27798 13268 27804 13280
rect 27856 13268 27862 13320
rect 28644 13317 28672 13348
rect 28920 13320 28948 13416
rect 29086 13336 29092 13388
rect 29144 13376 29150 13388
rect 30101 13379 30159 13385
rect 30101 13376 30113 13379
rect 29144 13348 30113 13376
rect 29144 13336 29150 13348
rect 30101 13345 30113 13348
rect 30147 13345 30159 13379
rect 30944 13376 30972 13416
rect 31662 13404 31668 13416
rect 31720 13404 31726 13456
rect 33594 13404 33600 13456
rect 33652 13444 33658 13456
rect 39114 13444 39120 13456
rect 33652 13416 39120 13444
rect 33652 13404 33658 13416
rect 39114 13404 39120 13416
rect 39172 13404 39178 13456
rect 43088 13444 43116 13472
rect 44358 13444 44364 13456
rect 43088 13416 43484 13444
rect 30944 13348 31064 13376
rect 30101 13339 30159 13345
rect 27985 13311 28043 13317
rect 27985 13277 27997 13311
rect 28031 13277 28043 13311
rect 27985 13271 28043 13277
rect 28629 13311 28687 13317
rect 28629 13277 28641 13311
rect 28675 13277 28687 13311
rect 28629 13271 28687 13277
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13277 28779 13311
rect 28902 13308 28908 13320
rect 28863 13280 28908 13308
rect 28721 13271 28779 13277
rect 24854 13240 24860 13252
rect 24815 13212 24860 13240
rect 24854 13200 24860 13212
rect 24912 13200 24918 13252
rect 26970 13240 26976 13252
rect 26931 13212 26976 13240
rect 26970 13200 26976 13212
rect 27028 13200 27034 13252
rect 24029 13175 24087 13181
rect 24029 13141 24041 13175
rect 24075 13172 24087 13175
rect 24486 13172 24492 13184
rect 24075 13144 24492 13172
rect 24075 13141 24087 13144
rect 24029 13135 24087 13141
rect 24486 13132 24492 13144
rect 24544 13132 24550 13184
rect 27706 13132 27712 13184
rect 27764 13172 27770 13184
rect 27893 13175 27951 13181
rect 27893 13172 27905 13175
rect 27764 13144 27905 13172
rect 27764 13132 27770 13144
rect 27893 13141 27905 13144
rect 27939 13141 27951 13175
rect 28000 13172 28028 13271
rect 28736 13240 28764 13271
rect 28902 13268 28908 13280
rect 28960 13268 28966 13320
rect 28994 13268 29000 13320
rect 29052 13308 29058 13320
rect 29181 13311 29239 13317
rect 29052 13280 29097 13308
rect 29052 13268 29058 13280
rect 29181 13277 29193 13311
rect 29227 13308 29239 13311
rect 29362 13308 29368 13320
rect 29227 13280 29368 13308
rect 29227 13277 29239 13280
rect 29181 13271 29239 13277
rect 29362 13268 29368 13280
rect 29420 13268 29426 13320
rect 29822 13268 29828 13320
rect 29880 13308 29886 13320
rect 29917 13311 29975 13317
rect 29917 13308 29929 13311
rect 29880 13280 29929 13308
rect 29880 13268 29886 13280
rect 29917 13277 29929 13280
rect 29963 13277 29975 13311
rect 29917 13271 29975 13277
rect 30653 13311 30711 13317
rect 30653 13277 30665 13311
rect 30699 13277 30711 13311
rect 30834 13308 30840 13320
rect 30795 13280 30840 13308
rect 30653 13271 30711 13277
rect 29733 13243 29791 13249
rect 29733 13240 29745 13243
rect 28736 13212 29745 13240
rect 29733 13209 29745 13212
rect 29779 13209 29791 13243
rect 30668 13240 30696 13271
rect 30834 13268 30840 13280
rect 30892 13268 30898 13320
rect 31036 13317 31064 13348
rect 33042 13336 33048 13388
rect 33100 13376 33106 13388
rect 34333 13379 34391 13385
rect 34333 13376 34345 13379
rect 33100 13348 34345 13376
rect 33100 13336 33106 13348
rect 34333 13345 34345 13348
rect 34379 13376 34391 13379
rect 34379 13348 35388 13376
rect 34379 13345 34391 13348
rect 34333 13339 34391 13345
rect 30929 13311 30987 13317
rect 30929 13277 30941 13311
rect 30975 13277 30987 13311
rect 30929 13271 30987 13277
rect 31021 13311 31079 13317
rect 31021 13277 31033 13311
rect 31067 13308 31079 13311
rect 31849 13311 31907 13317
rect 31849 13308 31861 13311
rect 31067 13280 31861 13308
rect 31067 13277 31079 13280
rect 31021 13271 31079 13277
rect 31849 13277 31861 13280
rect 31895 13308 31907 13311
rect 33226 13308 33232 13320
rect 31895 13280 33232 13308
rect 31895 13277 31907 13280
rect 31849 13271 31907 13277
rect 30742 13240 30748 13252
rect 30668 13212 30748 13240
rect 29733 13203 29791 13209
rect 30742 13200 30748 13212
rect 30800 13200 30806 13252
rect 30944 13240 30972 13271
rect 33226 13268 33232 13280
rect 33284 13308 33290 13320
rect 33870 13311 33928 13317
rect 33870 13308 33882 13311
rect 33284 13280 33882 13308
rect 33284 13268 33290 13280
rect 33870 13277 33882 13280
rect 33916 13308 33928 13311
rect 33962 13308 33968 13320
rect 33916 13280 33968 13308
rect 33916 13277 33928 13280
rect 33870 13271 33928 13277
rect 33962 13268 33968 13280
rect 34020 13268 34026 13320
rect 34238 13308 34244 13320
rect 34151 13280 34244 13308
rect 34238 13268 34244 13280
rect 34296 13308 34302 13320
rect 34296 13280 35296 13308
rect 34296 13268 34302 13280
rect 35158 13240 35164 13252
rect 30944 13212 35164 13240
rect 35158 13200 35164 13212
rect 35216 13200 35222 13252
rect 29178 13172 29184 13184
rect 28000 13144 29184 13172
rect 27893 13135 27951 13141
rect 29178 13132 29184 13144
rect 29236 13132 29242 13184
rect 33502 13132 33508 13184
rect 33560 13172 33566 13184
rect 33873 13175 33931 13181
rect 33873 13172 33885 13175
rect 33560 13144 33885 13172
rect 33560 13132 33566 13144
rect 33873 13141 33885 13144
rect 33919 13172 33931 13175
rect 34330 13172 34336 13184
rect 33919 13144 34336 13172
rect 33919 13141 33931 13144
rect 33873 13135 33931 13141
rect 34330 13132 34336 13144
rect 34388 13132 34394 13184
rect 34977 13175 35035 13181
rect 34977 13141 34989 13175
rect 35023 13172 35035 13175
rect 35268 13172 35296 13280
rect 35360 13240 35388 13348
rect 37182 13336 37188 13388
rect 37240 13376 37246 13388
rect 37369 13379 37427 13385
rect 37369 13376 37381 13379
rect 37240 13348 37381 13376
rect 37240 13336 37246 13348
rect 37369 13345 37381 13348
rect 37415 13345 37427 13379
rect 37369 13339 37427 13345
rect 37553 13379 37611 13385
rect 37553 13345 37565 13379
rect 37599 13376 37611 13379
rect 38654 13376 38660 13388
rect 37599 13348 38660 13376
rect 37599 13345 37611 13348
rect 37553 13339 37611 13345
rect 38654 13336 38660 13348
rect 38712 13336 38718 13388
rect 40402 13336 40408 13388
rect 40460 13376 40466 13388
rect 40497 13379 40555 13385
rect 40497 13376 40509 13379
rect 40460 13348 40509 13376
rect 40460 13336 40466 13348
rect 40497 13345 40509 13348
rect 40543 13345 40555 13379
rect 40497 13339 40555 13345
rect 40681 13379 40739 13385
rect 40681 13345 40693 13379
rect 40727 13376 40739 13379
rect 41230 13376 41236 13388
rect 40727 13348 41236 13376
rect 40727 13345 40739 13348
rect 40681 13339 40739 13345
rect 41230 13336 41236 13348
rect 41288 13336 41294 13388
rect 42521 13379 42579 13385
rect 42521 13345 42533 13379
rect 42567 13376 42579 13379
rect 43346 13376 43352 13388
rect 42567 13348 43352 13376
rect 42567 13345 42579 13348
rect 42521 13339 42579 13345
rect 43346 13336 43352 13348
rect 43404 13336 43410 13388
rect 35434 13268 35440 13320
rect 35492 13308 35498 13320
rect 35492 13280 35537 13308
rect 35492 13268 35498 13280
rect 36170 13268 36176 13320
rect 36228 13308 36234 13320
rect 37277 13311 37335 13317
rect 37277 13308 37289 13311
rect 36228 13280 37289 13308
rect 36228 13268 36234 13280
rect 37277 13277 37289 13280
rect 37323 13277 37335 13311
rect 37277 13271 37335 13277
rect 38013 13311 38071 13317
rect 38013 13277 38025 13311
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 38197 13311 38255 13317
rect 38197 13277 38209 13311
rect 38243 13308 38255 13311
rect 41966 13308 41972 13320
rect 38243 13280 38608 13308
rect 41927 13280 41972 13308
rect 38243 13277 38255 13280
rect 38197 13271 38255 13277
rect 36633 13243 36691 13249
rect 36633 13240 36645 13243
rect 35360 13212 36645 13240
rect 36633 13209 36645 13212
rect 36679 13240 36691 13243
rect 36722 13240 36728 13252
rect 36679 13212 36728 13240
rect 36679 13209 36691 13212
rect 36633 13203 36691 13209
rect 36722 13200 36728 13212
rect 36780 13200 36786 13252
rect 36814 13200 36820 13252
rect 36872 13240 36878 13252
rect 38028 13240 38056 13271
rect 36872 13212 38056 13240
rect 36872 13200 36878 13212
rect 38580 13184 38608 13280
rect 41966 13268 41972 13280
rect 42024 13268 42030 13320
rect 42337 13311 42395 13317
rect 42337 13277 42349 13311
rect 42383 13277 42395 13311
rect 42978 13308 42984 13320
rect 42939 13280 42984 13308
rect 42337 13271 42395 13277
rect 40218 13200 40224 13252
rect 40276 13240 40282 13252
rect 41233 13243 41291 13249
rect 41233 13240 41245 13243
rect 40276 13212 41245 13240
rect 40276 13200 40282 13212
rect 41233 13209 41245 13212
rect 41279 13209 41291 13243
rect 42352 13240 42380 13271
rect 42978 13268 42984 13280
rect 43036 13268 43042 13320
rect 43162 13308 43168 13320
rect 43123 13280 43168 13308
rect 43162 13268 43168 13280
rect 43220 13268 43226 13320
rect 43180 13240 43208 13268
rect 42352 13212 43208 13240
rect 43456 13240 43484 13416
rect 43640 13416 44364 13444
rect 43640 13317 43668 13416
rect 44358 13404 44364 13416
rect 44416 13404 44422 13456
rect 45922 13404 45928 13456
rect 45980 13404 45986 13456
rect 46014 13404 46020 13456
rect 46072 13404 46078 13456
rect 46216 13444 46244 13484
rect 46382 13472 46388 13484
rect 46440 13472 46446 13524
rect 47118 13472 47124 13524
rect 47176 13512 47182 13524
rect 47305 13515 47363 13521
rect 47305 13512 47317 13515
rect 47176 13484 47317 13512
rect 47176 13472 47182 13484
rect 47305 13481 47317 13484
rect 47351 13481 47363 13515
rect 47305 13475 47363 13481
rect 48038 13472 48044 13524
rect 48096 13512 48102 13524
rect 48498 13512 48504 13524
rect 48096 13484 48504 13512
rect 48096 13472 48102 13484
rect 48498 13472 48504 13484
rect 48556 13472 48562 13524
rect 48682 13512 48688 13524
rect 48643 13484 48688 13512
rect 48682 13472 48688 13484
rect 48740 13472 48746 13524
rect 50062 13512 50068 13524
rect 48884 13484 50068 13512
rect 47210 13444 47216 13456
rect 46216 13416 47216 13444
rect 47210 13404 47216 13416
rect 47268 13404 47274 13456
rect 48884 13444 48912 13484
rect 50062 13472 50068 13484
rect 50120 13512 50126 13524
rect 50430 13512 50436 13524
rect 50120 13484 50436 13512
rect 50120 13472 50126 13484
rect 50430 13472 50436 13484
rect 50488 13472 50494 13524
rect 50982 13472 50988 13524
rect 51040 13512 51046 13524
rect 51350 13512 51356 13524
rect 51040 13484 51356 13512
rect 51040 13472 51046 13484
rect 51350 13472 51356 13484
rect 51408 13472 51414 13524
rect 52178 13512 52184 13524
rect 52139 13484 52184 13512
rect 52178 13472 52184 13484
rect 52236 13472 52242 13524
rect 52822 13472 52828 13524
rect 52880 13512 52886 13524
rect 54386 13512 54392 13524
rect 52880 13484 54392 13512
rect 52880 13472 52886 13484
rect 54386 13472 54392 13484
rect 54444 13472 54450 13524
rect 54570 13472 54576 13524
rect 54628 13512 54634 13524
rect 54665 13515 54723 13521
rect 54665 13512 54677 13515
rect 54628 13484 54677 13512
rect 54628 13472 54634 13484
rect 54665 13481 54677 13484
rect 54711 13481 54723 13515
rect 56502 13512 56508 13524
rect 54665 13475 54723 13481
rect 55968 13484 56508 13512
rect 47504 13416 48912 13444
rect 43898 13336 43904 13388
rect 43956 13376 43962 13388
rect 43956 13348 44020 13376
rect 43956 13336 43962 13348
rect 43806 13317 43812 13320
rect 43625 13311 43683 13317
rect 43625 13277 43637 13311
rect 43671 13277 43683 13311
rect 43625 13271 43683 13277
rect 43773 13311 43812 13317
rect 43773 13277 43785 13311
rect 43773 13271 43812 13277
rect 43806 13268 43812 13271
rect 43864 13268 43870 13320
rect 43992 13317 44020 13348
rect 44542 13336 44548 13388
rect 44600 13376 44606 13388
rect 44600 13348 44956 13376
rect 44600 13336 44606 13348
rect 43992 13311 44051 13317
rect 43992 13277 44005 13311
rect 44039 13277 44051 13311
rect 43993 13271 44051 13277
rect 44131 13311 44189 13317
rect 44131 13277 44143 13311
rect 44177 13308 44189 13311
rect 44634 13308 44640 13320
rect 44177 13280 44640 13308
rect 44177 13277 44189 13280
rect 44131 13271 44189 13277
rect 44634 13268 44640 13280
rect 44692 13268 44698 13320
rect 44928 13308 44956 13348
rect 45370 13308 45376 13320
rect 44928 13280 45376 13308
rect 45370 13268 45376 13280
rect 45428 13308 45434 13320
rect 45940 13317 45968 13404
rect 46019 13317 46047 13404
rect 46382 13336 46388 13388
rect 46440 13376 46446 13388
rect 46750 13376 46756 13388
rect 46440 13348 46756 13376
rect 46440 13336 46446 13348
rect 46750 13336 46756 13348
rect 46808 13336 46814 13388
rect 47504 13317 47532 13416
rect 48958 13404 48964 13456
rect 49016 13444 49022 13456
rect 53653 13447 53711 13453
rect 53653 13444 53665 13447
rect 49016 13416 53665 13444
rect 49016 13404 49022 13416
rect 47946 13336 47952 13388
rect 48004 13376 48010 13388
rect 48498 13376 48504 13388
rect 48004 13348 48504 13376
rect 48004 13336 48010 13348
rect 48498 13336 48504 13348
rect 48556 13336 48562 13388
rect 45741 13311 45799 13317
rect 45741 13308 45753 13311
rect 45428 13280 45753 13308
rect 45428 13268 45434 13280
rect 45741 13277 45753 13280
rect 45787 13277 45799 13311
rect 45741 13271 45799 13277
rect 45904 13311 45968 13317
rect 45904 13277 45916 13311
rect 45950 13280 45968 13311
rect 46004 13311 46062 13317
rect 45950 13277 45962 13280
rect 45904 13271 45962 13277
rect 46004 13277 46016 13311
rect 46050 13277 46062 13311
rect 46004 13271 46062 13277
rect 46109 13311 46167 13317
rect 46109 13277 46121 13311
rect 46155 13277 46167 13311
rect 46109 13271 46167 13277
rect 47489 13311 47547 13317
rect 47489 13277 47501 13311
rect 47535 13277 47547 13311
rect 47489 13271 47547 13277
rect 47581 13311 47639 13317
rect 47581 13277 47593 13311
rect 47627 13277 47639 13311
rect 47581 13271 47639 13277
rect 47765 13311 47823 13317
rect 47765 13277 47777 13311
rect 47811 13277 47823 13311
rect 47765 13271 47823 13277
rect 47857 13311 47915 13317
rect 47857 13277 47869 13311
rect 47903 13308 47915 13311
rect 48130 13308 48136 13320
rect 47903 13280 48136 13308
rect 47903 13277 47915 13280
rect 47857 13271 47915 13277
rect 43901 13243 43959 13249
rect 43901 13240 43913 13243
rect 43456 13212 43913 13240
rect 41233 13203 41291 13209
rect 38010 13172 38016 13184
rect 35023 13144 38016 13172
rect 35023 13141 35035 13144
rect 34977 13135 35035 13141
rect 38010 13132 38016 13144
rect 38068 13132 38074 13184
rect 38105 13175 38163 13181
rect 38105 13141 38117 13175
rect 38151 13172 38163 13175
rect 38286 13172 38292 13184
rect 38151 13144 38292 13172
rect 38151 13141 38163 13144
rect 38105 13135 38163 13141
rect 38286 13132 38292 13144
rect 38344 13132 38350 13184
rect 38562 13132 38568 13184
rect 38620 13172 38626 13184
rect 38657 13175 38715 13181
rect 38657 13172 38669 13175
rect 38620 13144 38669 13172
rect 38620 13132 38626 13144
rect 38657 13141 38669 13144
rect 38703 13141 38715 13175
rect 38657 13135 38715 13141
rect 40405 13175 40463 13181
rect 40405 13141 40417 13175
rect 40451 13172 40463 13175
rect 40770 13172 40776 13184
rect 40451 13144 40776 13172
rect 40451 13141 40463 13144
rect 40405 13135 40463 13141
rect 40770 13132 40776 13144
rect 40828 13132 40834 13184
rect 42334 13172 42340 13184
rect 42295 13144 42340 13172
rect 42334 13132 42340 13144
rect 42392 13132 42398 13184
rect 43180 13172 43208 13212
rect 43901 13209 43913 13212
rect 43947 13209 43959 13243
rect 43901 13203 43959 13209
rect 45646 13200 45652 13252
rect 45704 13240 45710 13252
rect 45704 13212 46047 13240
rect 45704 13200 45710 13212
rect 45186 13172 45192 13184
rect 43180 13144 45192 13172
rect 45186 13132 45192 13144
rect 45244 13132 45250 13184
rect 46019 13172 46047 13212
rect 46124 13172 46152 13271
rect 47026 13200 47032 13252
rect 47084 13240 47090 13252
rect 47596 13240 47624 13271
rect 47084 13212 47624 13240
rect 47780 13240 47808 13271
rect 48130 13268 48136 13280
rect 48188 13268 48194 13320
rect 48222 13268 48228 13320
rect 48280 13308 48286 13320
rect 49620 13317 49648 13416
rect 53653 13413 53665 13416
rect 53699 13444 53711 13447
rect 54202 13444 54208 13456
rect 53699 13416 54208 13444
rect 53699 13413 53711 13416
rect 53653 13407 53711 13413
rect 54202 13404 54208 13416
rect 54260 13404 54266 13456
rect 54481 13447 54539 13453
rect 54481 13413 54493 13447
rect 54527 13444 54539 13447
rect 55122 13444 55128 13456
rect 54527 13416 55128 13444
rect 54527 13413 54539 13416
rect 54481 13407 54539 13413
rect 49694 13336 49700 13388
rect 49752 13376 49758 13388
rect 51350 13376 51356 13388
rect 49752 13348 51356 13376
rect 49752 13336 49758 13348
rect 49605 13311 49663 13317
rect 48280 13280 49464 13308
rect 48280 13268 48286 13280
rect 48038 13240 48044 13252
rect 47780 13212 48044 13240
rect 47084 13200 47090 13212
rect 48038 13200 48044 13212
rect 48096 13200 48102 13252
rect 48317 13243 48375 13249
rect 48317 13209 48329 13243
rect 48363 13209 48375 13243
rect 48317 13203 48375 13209
rect 46019 13144 46152 13172
rect 46198 13132 46204 13184
rect 46256 13172 46262 13184
rect 48332 13172 48360 13203
rect 48498 13200 48504 13252
rect 48556 13240 48562 13252
rect 48682 13240 48688 13252
rect 48556 13212 48688 13240
rect 48556 13200 48562 13212
rect 48682 13200 48688 13212
rect 48740 13200 48746 13252
rect 49436 13181 49464 13280
rect 49605 13277 49617 13311
rect 49651 13277 49663 13311
rect 49605 13271 49663 13277
rect 49786 13268 49792 13320
rect 49844 13308 49850 13320
rect 50448 13317 50476 13348
rect 51350 13336 51356 13348
rect 51408 13336 51414 13388
rect 51810 13376 51816 13388
rect 51460 13348 51816 13376
rect 50341 13311 50399 13317
rect 50341 13308 50353 13311
rect 49844 13280 50353 13308
rect 49844 13268 49850 13280
rect 50341 13277 50353 13280
rect 50387 13277 50399 13311
rect 50341 13271 50399 13277
rect 50433 13311 50491 13317
rect 50433 13277 50445 13311
rect 50479 13277 50491 13311
rect 50433 13271 50491 13277
rect 50617 13311 50675 13317
rect 50617 13277 50629 13311
rect 50663 13308 50675 13311
rect 50706 13308 50712 13320
rect 50663 13280 50712 13308
rect 50663 13277 50675 13280
rect 50617 13271 50675 13277
rect 50706 13268 50712 13280
rect 50764 13308 50770 13320
rect 51460 13317 51488 13348
rect 51810 13336 51816 13348
rect 51868 13336 51874 13388
rect 52638 13336 52644 13388
rect 52696 13376 52702 13388
rect 53742 13376 53748 13388
rect 52696 13348 53748 13376
rect 52696 13336 52702 13348
rect 53742 13336 53748 13348
rect 53800 13336 53806 13388
rect 51261 13311 51319 13317
rect 51261 13308 51273 13311
rect 50764 13280 51273 13308
rect 50764 13268 50770 13280
rect 51261 13277 51273 13280
rect 51307 13277 51319 13311
rect 51261 13271 51319 13277
rect 51445 13311 51503 13317
rect 51445 13277 51457 13311
rect 51491 13277 51503 13311
rect 51445 13271 51503 13277
rect 51721 13311 51779 13317
rect 51721 13277 51733 13311
rect 51767 13277 51779 13311
rect 51721 13271 51779 13277
rect 49694 13200 49700 13252
rect 49752 13240 49758 13252
rect 50801 13243 50859 13249
rect 50801 13240 50813 13243
rect 49752 13212 50813 13240
rect 49752 13200 49758 13212
rect 50801 13209 50813 13212
rect 50847 13209 50859 13243
rect 51736 13240 51764 13271
rect 52454 13268 52460 13320
rect 52512 13308 52518 13320
rect 53190 13308 53196 13320
rect 52512 13280 53196 13308
rect 52512 13268 52518 13280
rect 53190 13268 53196 13280
rect 53248 13308 53254 13320
rect 53466 13308 53472 13320
rect 53248 13280 53472 13308
rect 53248 13268 53254 13280
rect 53466 13268 53472 13280
rect 53524 13268 53530 13320
rect 53561 13311 53619 13317
rect 53561 13277 53573 13311
rect 53607 13308 53619 13311
rect 54496 13308 54524 13407
rect 55122 13404 55128 13416
rect 55180 13404 55186 13456
rect 55493 13447 55551 13453
rect 55493 13413 55505 13447
rect 55539 13444 55551 13447
rect 55582 13444 55588 13456
rect 55539 13416 55588 13444
rect 55539 13413 55551 13416
rect 55493 13407 55551 13413
rect 55582 13404 55588 13416
rect 55640 13404 55646 13456
rect 55968 13376 55996 13484
rect 56502 13472 56508 13484
rect 56560 13472 56566 13524
rect 56594 13472 56600 13524
rect 56652 13512 56658 13524
rect 56652 13484 56697 13512
rect 56652 13472 56658 13484
rect 56410 13444 56416 13456
rect 55876 13348 55996 13376
rect 56060 13416 56416 13444
rect 55876 13317 55904 13348
rect 53607 13280 54524 13308
rect 55861 13311 55919 13317
rect 55768 13289 55826 13295
rect 53607 13277 53619 13280
rect 53561 13271 53619 13277
rect 55768 13255 55780 13289
rect 55814 13286 55826 13289
rect 55814 13255 55828 13286
rect 55861 13277 55873 13311
rect 55907 13277 55919 13311
rect 55861 13271 55919 13277
rect 55953 13311 56011 13317
rect 55953 13277 55965 13311
rect 55999 13308 56011 13311
rect 56060 13308 56088 13416
rect 56410 13404 56416 13416
rect 56468 13404 56474 13456
rect 55999 13280 56088 13308
rect 56137 13311 56195 13317
rect 55999 13277 56011 13280
rect 55953 13271 56011 13277
rect 56137 13277 56149 13311
rect 56183 13308 56195 13311
rect 56226 13308 56232 13320
rect 56183 13280 56232 13308
rect 56183 13277 56195 13280
rect 56137 13271 56195 13277
rect 56226 13268 56232 13280
rect 56284 13268 56290 13320
rect 57974 13268 57980 13320
rect 58032 13308 58038 13320
rect 58069 13311 58127 13317
rect 58069 13308 58081 13311
rect 58032 13280 58081 13308
rect 58032 13268 58038 13280
rect 58069 13277 58081 13280
rect 58115 13308 58127 13311
rect 58434 13308 58440 13320
rect 58115 13280 58440 13308
rect 58115 13277 58127 13280
rect 58069 13271 58127 13277
rect 58434 13268 58440 13280
rect 58492 13268 58498 13320
rect 51736 13212 54156 13240
rect 50801 13203 50859 13209
rect 46256 13144 48360 13172
rect 49421 13175 49479 13181
rect 46256 13132 46262 13144
rect 49421 13141 49433 13175
rect 49467 13141 49479 13175
rect 49421 13135 49479 13141
rect 49602 13132 49608 13184
rect 49660 13172 49666 13184
rect 51166 13172 51172 13184
rect 49660 13144 51172 13172
rect 49660 13132 49666 13144
rect 51166 13132 51172 13144
rect 51224 13172 51230 13184
rect 51442 13172 51448 13184
rect 51224 13144 51448 13172
rect 51224 13132 51230 13144
rect 51442 13132 51448 13144
rect 51500 13172 51506 13184
rect 51629 13175 51687 13181
rect 51629 13172 51641 13175
rect 51500 13144 51641 13172
rect 51500 13132 51506 13144
rect 51629 13141 51641 13144
rect 51675 13141 51687 13175
rect 51629 13135 51687 13141
rect 52546 13132 52552 13184
rect 52604 13172 52610 13184
rect 52733 13175 52791 13181
rect 52733 13172 52745 13175
rect 52604 13144 52745 13172
rect 52604 13132 52610 13144
rect 52733 13141 52745 13144
rect 52779 13141 52791 13175
rect 52733 13135 52791 13141
rect 53190 13132 53196 13184
rect 53248 13172 53254 13184
rect 53650 13172 53656 13184
rect 53248 13144 53656 13172
rect 53248 13132 53254 13144
rect 53650 13132 53656 13144
rect 53708 13132 53714 13184
rect 54128 13172 54156 13212
rect 54202 13200 54208 13252
rect 54260 13240 54266 13252
rect 55768 13249 55828 13255
rect 55800 13240 55828 13249
rect 56042 13240 56048 13252
rect 54260 13212 54305 13240
rect 55800 13212 56048 13240
rect 54260 13200 54266 13212
rect 56042 13200 56048 13212
rect 56100 13200 56106 13252
rect 55858 13172 55864 13184
rect 54128 13144 55864 13172
rect 55858 13132 55864 13144
rect 55916 13132 55922 13184
rect 56226 13132 56232 13184
rect 56284 13172 56290 13184
rect 57149 13175 57207 13181
rect 57149 13172 57161 13175
rect 56284 13144 57161 13172
rect 56284 13132 56290 13144
rect 57149 13141 57161 13144
rect 57195 13141 57207 13175
rect 58250 13172 58256 13184
rect 58211 13144 58256 13172
rect 57149 13135 57207 13141
rect 58250 13132 58256 13144
rect 58308 13132 58314 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 25866 12968 25872 12980
rect 25827 12940 25872 12968
rect 25866 12928 25872 12940
rect 25924 12928 25930 12980
rect 26142 12928 26148 12980
rect 26200 12968 26206 12980
rect 27890 12968 27896 12980
rect 26200 12940 27896 12968
rect 26200 12928 26206 12940
rect 27890 12928 27896 12940
rect 27948 12968 27954 12980
rect 28445 12971 28503 12977
rect 28445 12968 28457 12971
rect 27948 12940 28457 12968
rect 27948 12928 27954 12940
rect 28445 12937 28457 12940
rect 28491 12968 28503 12971
rect 28902 12968 28908 12980
rect 28491 12940 28908 12968
rect 28491 12937 28503 12940
rect 28445 12931 28503 12937
rect 28902 12928 28908 12940
rect 28960 12928 28966 12980
rect 29089 12971 29147 12977
rect 29089 12937 29101 12971
rect 29135 12968 29147 12971
rect 29178 12968 29184 12980
rect 29135 12940 29184 12968
rect 29135 12937 29147 12940
rect 29089 12931 29147 12937
rect 29178 12928 29184 12940
rect 29236 12928 29242 12980
rect 31297 12971 31355 12977
rect 31297 12937 31309 12971
rect 31343 12968 31355 12971
rect 31846 12968 31852 12980
rect 31343 12940 31852 12968
rect 31343 12937 31355 12940
rect 31297 12931 31355 12937
rect 31846 12928 31852 12940
rect 31904 12928 31910 12980
rect 33321 12971 33379 12977
rect 33321 12937 33333 12971
rect 33367 12968 33379 12971
rect 33410 12968 33416 12980
rect 33367 12940 33416 12968
rect 33367 12937 33379 12940
rect 33321 12931 33379 12937
rect 33410 12928 33416 12940
rect 33468 12928 33474 12980
rect 34238 12968 34244 12980
rect 34199 12940 34244 12968
rect 34238 12928 34244 12940
rect 34296 12928 34302 12980
rect 34514 12928 34520 12980
rect 34572 12968 34578 12980
rect 35342 12968 35348 12980
rect 34572 12940 35348 12968
rect 34572 12928 34578 12940
rect 35342 12928 35348 12940
rect 35400 12928 35406 12980
rect 35713 12971 35771 12977
rect 35713 12937 35725 12971
rect 35759 12968 35771 12971
rect 35894 12968 35900 12980
rect 35759 12940 35900 12968
rect 35759 12937 35771 12940
rect 35713 12931 35771 12937
rect 35894 12928 35900 12940
rect 35952 12928 35958 12980
rect 36173 12971 36231 12977
rect 36173 12937 36185 12971
rect 36219 12968 36231 12971
rect 36446 12968 36452 12980
rect 36219 12940 36452 12968
rect 36219 12937 36231 12940
rect 36173 12931 36231 12937
rect 36446 12928 36452 12940
rect 36504 12928 36510 12980
rect 37918 12928 37924 12980
rect 37976 12968 37982 12980
rect 40218 12968 40224 12980
rect 37976 12940 40224 12968
rect 37976 12928 37982 12940
rect 40218 12928 40224 12940
rect 40276 12928 40282 12980
rect 40494 12928 40500 12980
rect 40552 12968 40558 12980
rect 40957 12971 41015 12977
rect 40957 12968 40969 12971
rect 40552 12940 40969 12968
rect 40552 12928 40558 12940
rect 40957 12937 40969 12940
rect 41003 12937 41015 12971
rect 42702 12968 42708 12980
rect 42663 12940 42708 12968
rect 40957 12931 41015 12937
rect 42702 12928 42708 12940
rect 42760 12928 42766 12980
rect 43073 12971 43131 12977
rect 43073 12937 43085 12971
rect 43119 12968 43131 12971
rect 44542 12968 44548 12980
rect 43119 12940 44548 12968
rect 43119 12937 43131 12940
rect 43073 12931 43131 12937
rect 24949 12903 25007 12909
rect 24949 12869 24961 12903
rect 24995 12900 25007 12903
rect 28074 12900 28080 12912
rect 24995 12872 26280 12900
rect 24995 12869 25007 12872
rect 24949 12863 25007 12869
rect 23753 12835 23811 12841
rect 23753 12832 23765 12835
rect 6886 12804 23765 12832
rect 1854 12588 1860 12640
rect 1912 12628 1918 12640
rect 6886 12628 6914 12804
rect 23753 12801 23765 12804
rect 23799 12832 23811 12835
rect 24302 12832 24308 12844
rect 23799 12804 24308 12832
rect 23799 12801 23811 12804
rect 23753 12795 23811 12801
rect 24302 12792 24308 12804
rect 24360 12792 24366 12844
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 24854 12832 24860 12844
rect 24443 12804 24860 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 24854 12792 24860 12804
rect 24912 12832 24918 12844
rect 25133 12835 25191 12841
rect 25133 12832 25145 12835
rect 24912 12804 25145 12832
rect 24912 12792 24918 12804
rect 25133 12801 25145 12804
rect 25179 12801 25191 12835
rect 25133 12795 25191 12801
rect 25317 12835 25375 12841
rect 25317 12801 25329 12835
rect 25363 12832 25375 12835
rect 25958 12832 25964 12844
rect 25363 12804 25964 12832
rect 25363 12801 25375 12804
rect 25317 12795 25375 12801
rect 24486 12724 24492 12776
rect 24544 12764 24550 12776
rect 25332 12764 25360 12795
rect 25958 12792 25964 12804
rect 26016 12792 26022 12844
rect 26050 12792 26056 12844
rect 26108 12832 26114 12844
rect 26252 12841 26280 12872
rect 27816 12872 28080 12900
rect 26237 12835 26295 12841
rect 26108 12804 26153 12832
rect 26108 12792 26114 12804
rect 26237 12801 26249 12835
rect 26283 12801 26295 12835
rect 26237 12795 26295 12801
rect 26418 12792 26424 12844
rect 26476 12832 26482 12844
rect 26513 12835 26571 12841
rect 26513 12832 26525 12835
rect 26476 12804 26525 12832
rect 26476 12792 26482 12804
rect 26513 12801 26525 12804
rect 26559 12801 26571 12835
rect 27154 12832 27160 12844
rect 27115 12804 27160 12832
rect 26513 12795 26571 12801
rect 27154 12792 27160 12804
rect 27212 12792 27218 12844
rect 27430 12832 27436 12844
rect 27391 12804 27436 12832
rect 27430 12792 27436 12804
rect 27488 12792 27494 12844
rect 27706 12832 27712 12844
rect 27667 12804 27712 12832
rect 27706 12792 27712 12804
rect 27764 12792 27770 12844
rect 24544 12736 25360 12764
rect 25409 12767 25467 12773
rect 24544 12724 24550 12736
rect 25409 12733 25421 12767
rect 25455 12733 25467 12767
rect 25409 12727 25467 12733
rect 26329 12767 26387 12773
rect 26329 12733 26341 12767
rect 26375 12764 26387 12767
rect 27617 12767 27675 12773
rect 26375 12736 27384 12764
rect 26375 12733 26387 12736
rect 26329 12727 26387 12733
rect 1912 12600 6914 12628
rect 25424 12628 25452 12727
rect 27356 12708 27384 12736
rect 27617 12733 27629 12767
rect 27663 12764 27675 12767
rect 27816 12764 27844 12872
rect 28074 12860 28080 12872
rect 28132 12860 28138 12912
rect 34256 12900 34284 12928
rect 39390 12900 39396 12912
rect 29196 12872 33640 12900
rect 27893 12835 27951 12841
rect 27893 12801 27905 12835
rect 27939 12832 27951 12835
rect 28166 12832 28172 12844
rect 27939 12804 28172 12832
rect 27939 12801 27951 12804
rect 27893 12795 27951 12801
rect 28166 12792 28172 12804
rect 28224 12792 28230 12844
rect 28997 12835 29055 12841
rect 28997 12801 29009 12835
rect 29043 12832 29055 12835
rect 29086 12832 29092 12844
rect 29043 12804 29092 12832
rect 29043 12801 29055 12804
rect 28997 12795 29055 12801
rect 29086 12792 29092 12804
rect 29144 12792 29150 12844
rect 29196 12841 29224 12872
rect 33612 12844 33640 12872
rect 34164 12872 34284 12900
rect 35268 12872 35848 12900
rect 29181 12835 29239 12841
rect 29181 12801 29193 12835
rect 29227 12801 29239 12835
rect 29181 12795 29239 12801
rect 29454 12792 29460 12844
rect 29512 12832 29518 12844
rect 29641 12835 29699 12841
rect 29641 12832 29653 12835
rect 29512 12804 29653 12832
rect 29512 12792 29518 12804
rect 29641 12801 29653 12804
rect 29687 12801 29699 12835
rect 29822 12832 29828 12844
rect 29783 12804 29828 12832
rect 29641 12795 29699 12801
rect 29822 12792 29828 12804
rect 29880 12792 29886 12844
rect 30098 12792 30104 12844
rect 30156 12832 30162 12844
rect 31113 12835 31171 12841
rect 31113 12832 31125 12835
rect 30156 12804 31125 12832
rect 30156 12792 30162 12804
rect 31113 12801 31125 12804
rect 31159 12801 31171 12835
rect 32677 12835 32735 12841
rect 32677 12832 32689 12835
rect 31113 12795 31171 12801
rect 31726 12804 32689 12832
rect 27663 12736 27844 12764
rect 27663 12733 27675 12736
rect 27617 12727 27675 12733
rect 27982 12724 27988 12776
rect 28040 12764 28046 12776
rect 28040 12736 28856 12764
rect 28040 12724 28046 12736
rect 26145 12699 26203 12705
rect 26145 12665 26157 12699
rect 26191 12696 26203 12699
rect 27246 12696 27252 12708
rect 26191 12668 27252 12696
rect 26191 12665 26203 12668
rect 26145 12659 26203 12665
rect 27246 12656 27252 12668
rect 27304 12656 27310 12708
rect 27338 12656 27344 12708
rect 27396 12696 27402 12708
rect 28828 12696 28856 12736
rect 29546 12724 29552 12776
rect 29604 12764 29610 12776
rect 30837 12767 30895 12773
rect 30837 12764 30849 12767
rect 29604 12736 30849 12764
rect 29604 12724 29610 12736
rect 30837 12733 30849 12736
rect 30883 12764 30895 12767
rect 31726 12764 31754 12804
rect 32677 12801 32689 12804
rect 32723 12801 32735 12835
rect 32677 12795 32735 12801
rect 33505 12835 33563 12841
rect 33505 12801 33517 12835
rect 33551 12801 33563 12835
rect 33505 12795 33563 12801
rect 32490 12764 32496 12776
rect 30883 12736 31754 12764
rect 32451 12736 32496 12764
rect 30883 12733 30895 12736
rect 30837 12727 30895 12733
rect 32490 12724 32496 12736
rect 32548 12724 32554 12776
rect 32582 12724 32588 12776
rect 32640 12764 32646 12776
rect 32769 12767 32827 12773
rect 32640 12736 32685 12764
rect 32640 12724 32646 12736
rect 32769 12733 32781 12767
rect 32815 12764 32827 12767
rect 33520 12764 33548 12795
rect 33594 12792 33600 12844
rect 33652 12832 33658 12844
rect 33781 12835 33839 12841
rect 33652 12804 33697 12832
rect 33652 12792 33658 12804
rect 33781 12801 33793 12835
rect 33827 12832 33839 12835
rect 33962 12832 33968 12844
rect 33827 12804 33968 12832
rect 33827 12801 33839 12804
rect 33781 12795 33839 12801
rect 33962 12792 33968 12804
rect 34020 12792 34026 12844
rect 34164 12764 34192 12872
rect 34330 12792 34336 12844
rect 34388 12832 34394 12844
rect 34974 12832 34980 12844
rect 34388 12804 34980 12832
rect 34388 12792 34394 12804
rect 34974 12792 34980 12804
rect 35032 12792 35038 12844
rect 35158 12832 35164 12844
rect 35119 12804 35164 12832
rect 35158 12792 35164 12804
rect 35216 12832 35222 12844
rect 35268 12832 35296 12872
rect 35216 12804 35296 12832
rect 35529 12835 35587 12841
rect 35216 12792 35222 12804
rect 35529 12801 35541 12835
rect 35575 12832 35587 12835
rect 35710 12832 35716 12844
rect 35575 12804 35716 12832
rect 35575 12801 35587 12804
rect 35529 12795 35587 12801
rect 35710 12792 35716 12804
rect 35768 12792 35774 12844
rect 32815 12736 33456 12764
rect 33520 12736 34192 12764
rect 35253 12767 35311 12773
rect 32815 12733 32827 12736
rect 32769 12727 32827 12733
rect 32309 12699 32367 12705
rect 32309 12696 32321 12699
rect 27396 12668 28764 12696
rect 28828 12668 32321 12696
rect 27396 12656 27402 12668
rect 28736 12640 28764 12668
rect 32309 12665 32321 12668
rect 32355 12665 32367 12699
rect 32600 12696 32628 12724
rect 32858 12696 32864 12708
rect 32600 12668 32864 12696
rect 32309 12659 32367 12665
rect 32858 12656 32864 12668
rect 32916 12656 32922 12708
rect 33428 12696 33456 12736
rect 35253 12733 35265 12767
rect 35299 12733 35311 12767
rect 35253 12727 35311 12733
rect 35268 12696 35296 12727
rect 35342 12724 35348 12776
rect 35400 12764 35406 12776
rect 35820 12764 35848 12872
rect 38120 12872 39396 12900
rect 35894 12792 35900 12844
rect 35952 12832 35958 12844
rect 36078 12832 36084 12844
rect 35952 12804 36084 12832
rect 35952 12792 35958 12804
rect 36078 12792 36084 12804
rect 36136 12792 36142 12844
rect 36262 12792 36268 12844
rect 36320 12832 36326 12844
rect 36357 12835 36415 12841
rect 36357 12832 36369 12835
rect 36320 12804 36369 12832
rect 36320 12792 36326 12804
rect 36357 12801 36369 12804
rect 36403 12801 36415 12835
rect 36538 12832 36544 12844
rect 36499 12804 36544 12832
rect 36357 12795 36415 12801
rect 36538 12792 36544 12804
rect 36596 12792 36602 12844
rect 36630 12792 36636 12844
rect 36688 12832 36694 12844
rect 36688 12804 36733 12832
rect 36688 12792 36694 12804
rect 37182 12792 37188 12844
rect 37240 12832 37246 12844
rect 37553 12835 37611 12841
rect 37553 12832 37565 12835
rect 37240 12804 37565 12832
rect 37240 12792 37246 12804
rect 37553 12801 37565 12804
rect 37599 12832 37611 12835
rect 38013 12835 38071 12841
rect 38013 12832 38025 12835
rect 37599 12804 38025 12832
rect 37599 12801 37611 12804
rect 37553 12795 37611 12801
rect 38013 12801 38025 12804
rect 38059 12832 38071 12835
rect 38120 12832 38148 12872
rect 39390 12860 39396 12872
rect 39448 12860 39454 12912
rect 42610 12860 42616 12912
rect 42668 12900 42674 12912
rect 43088 12900 43116 12931
rect 44542 12928 44548 12940
rect 44600 12928 44606 12980
rect 44910 12928 44916 12980
rect 44968 12968 44974 12980
rect 45189 12971 45247 12977
rect 45189 12968 45201 12971
rect 44968 12940 45201 12968
rect 44968 12928 44974 12940
rect 45189 12937 45201 12940
rect 45235 12937 45247 12971
rect 45189 12931 45247 12937
rect 45922 12928 45928 12980
rect 45980 12968 45986 12980
rect 46293 12971 46351 12977
rect 46293 12968 46305 12971
rect 45980 12940 46305 12968
rect 45980 12928 45986 12940
rect 46293 12937 46305 12940
rect 46339 12937 46351 12971
rect 46293 12931 46351 12937
rect 47302 12928 47308 12980
rect 47360 12968 47366 12980
rect 47857 12971 47915 12977
rect 47857 12968 47869 12971
rect 47360 12940 47869 12968
rect 47360 12928 47366 12940
rect 47857 12937 47869 12940
rect 47903 12937 47915 12971
rect 49602 12968 49608 12980
rect 47857 12931 47915 12937
rect 49252 12940 49608 12968
rect 42668 12872 43116 12900
rect 43717 12903 43775 12909
rect 42668 12860 42674 12872
rect 43717 12869 43729 12903
rect 43763 12900 43775 12903
rect 43898 12900 43904 12912
rect 43763 12872 43904 12900
rect 43763 12869 43775 12872
rect 43717 12863 43775 12869
rect 43898 12860 43904 12872
rect 43956 12860 43962 12912
rect 44361 12903 44419 12909
rect 44361 12869 44373 12903
rect 44407 12900 44419 12903
rect 44634 12900 44640 12912
rect 44407 12872 44640 12900
rect 44407 12869 44419 12872
rect 44361 12863 44419 12869
rect 44634 12860 44640 12872
rect 44692 12860 44698 12912
rect 46014 12860 46020 12912
rect 46072 12900 46078 12912
rect 48222 12900 48228 12912
rect 46072 12872 48228 12900
rect 46072 12860 46078 12872
rect 48222 12860 48228 12872
rect 48280 12860 48286 12912
rect 48406 12860 48412 12912
rect 48464 12900 48470 12912
rect 49252 12900 49280 12940
rect 49602 12928 49608 12940
rect 49660 12928 49666 12980
rect 49878 12928 49884 12980
rect 49936 12968 49942 12980
rect 50525 12971 50583 12977
rect 50525 12968 50537 12971
rect 49936 12940 50537 12968
rect 49936 12928 49942 12940
rect 50525 12937 50537 12940
rect 50571 12937 50583 12971
rect 53834 12968 53840 12980
rect 50525 12931 50583 12937
rect 51046 12940 53840 12968
rect 48464 12872 49280 12900
rect 49329 12903 49387 12909
rect 48464 12860 48470 12872
rect 38059 12804 38148 12832
rect 38197 12835 38255 12841
rect 38059 12801 38071 12804
rect 38013 12795 38071 12801
rect 38197 12801 38209 12835
rect 38243 12832 38255 12835
rect 38286 12832 38292 12844
rect 38243 12804 38292 12832
rect 38243 12801 38255 12804
rect 38197 12795 38255 12801
rect 38286 12792 38292 12804
rect 38344 12832 38350 12844
rect 38749 12835 38807 12841
rect 38749 12832 38761 12835
rect 38344 12804 38761 12832
rect 38344 12792 38350 12804
rect 38749 12801 38761 12804
rect 38795 12801 38807 12835
rect 38749 12795 38807 12801
rect 39025 12835 39083 12841
rect 39025 12801 39037 12835
rect 39071 12832 39083 12835
rect 39206 12832 39212 12844
rect 39071 12804 39212 12832
rect 39071 12801 39083 12804
rect 39025 12795 39083 12801
rect 35400 12736 35445 12764
rect 35820 12736 36492 12764
rect 35400 12724 35406 12736
rect 36078 12696 36084 12708
rect 33428 12668 35204 12696
rect 35268 12668 36084 12696
rect 26786 12628 26792 12640
rect 25424 12600 26792 12628
rect 1912 12588 1918 12600
rect 26786 12588 26792 12600
rect 26844 12588 26850 12640
rect 28718 12588 28724 12640
rect 28776 12628 28782 12640
rect 29733 12631 29791 12637
rect 29733 12628 29745 12631
rect 28776 12600 29745 12628
rect 28776 12588 28782 12600
rect 29733 12597 29745 12600
rect 29779 12597 29791 12631
rect 29733 12591 29791 12597
rect 30374 12588 30380 12640
rect 30432 12628 30438 12640
rect 30742 12628 30748 12640
rect 30432 12600 30748 12628
rect 30432 12588 30438 12600
rect 30742 12588 30748 12600
rect 30800 12588 30806 12640
rect 30929 12631 30987 12637
rect 30929 12597 30941 12631
rect 30975 12628 30987 12631
rect 31018 12628 31024 12640
rect 30975 12600 31024 12628
rect 30975 12597 30987 12600
rect 30929 12591 30987 12597
rect 31018 12588 31024 12600
rect 31076 12588 31082 12640
rect 33781 12631 33839 12637
rect 33781 12597 33793 12631
rect 33827 12628 33839 12631
rect 34146 12628 34152 12640
rect 33827 12600 34152 12628
rect 33827 12597 33839 12600
rect 33781 12591 33839 12597
rect 34146 12588 34152 12600
rect 34204 12588 34210 12640
rect 35176 12628 35204 12668
rect 36078 12656 36084 12668
rect 36136 12656 36142 12708
rect 36464 12696 36492 12736
rect 36998 12724 37004 12776
rect 37056 12764 37062 12776
rect 38930 12764 38936 12776
rect 37056 12736 38792 12764
rect 38891 12736 38936 12764
rect 37056 12724 37062 12736
rect 38197 12699 38255 12705
rect 38197 12696 38209 12699
rect 36464 12668 38209 12696
rect 38197 12665 38209 12668
rect 38243 12665 38255 12699
rect 38764 12696 38792 12736
rect 38930 12724 38936 12736
rect 38988 12724 38994 12776
rect 39040 12696 39068 12795
rect 39206 12792 39212 12804
rect 39264 12792 39270 12844
rect 41785 12835 41843 12841
rect 41785 12801 41797 12835
rect 41831 12801 41843 12835
rect 42886 12832 42892 12844
rect 42847 12804 42892 12832
rect 41785 12795 41843 12801
rect 40497 12767 40555 12773
rect 40497 12733 40509 12767
rect 40543 12764 40555 12767
rect 40678 12764 40684 12776
rect 40543 12736 40684 12764
rect 40543 12733 40555 12736
rect 40497 12727 40555 12733
rect 40678 12724 40684 12736
rect 40736 12724 40742 12776
rect 41800 12764 41828 12795
rect 42886 12792 42892 12804
rect 42944 12832 42950 12844
rect 43070 12832 43076 12844
rect 42944 12804 43076 12832
rect 42944 12792 42950 12804
rect 43070 12792 43076 12804
rect 43128 12792 43134 12844
rect 43165 12835 43223 12841
rect 43165 12801 43177 12835
rect 43211 12832 43223 12835
rect 43254 12832 43260 12844
rect 43211 12804 43260 12832
rect 43211 12801 43223 12804
rect 43165 12795 43223 12801
rect 43254 12792 43260 12804
rect 43312 12792 43318 12844
rect 43622 12792 43628 12844
rect 43680 12832 43686 12844
rect 43809 12835 43867 12841
rect 43809 12832 43821 12835
rect 43680 12804 43821 12832
rect 43680 12792 43686 12804
rect 43809 12801 43821 12804
rect 43855 12801 43867 12835
rect 43809 12795 43867 12801
rect 45370 12792 45376 12844
rect 45428 12832 45434 12844
rect 45741 12835 45799 12841
rect 45741 12832 45753 12835
rect 45428 12804 45753 12832
rect 45428 12792 45434 12804
rect 45741 12801 45753 12804
rect 45787 12832 45799 12835
rect 46937 12835 46995 12841
rect 46937 12832 46949 12835
rect 45787 12804 46949 12832
rect 45787 12801 45799 12804
rect 45741 12795 45799 12801
rect 46937 12801 46949 12804
rect 46983 12801 46995 12835
rect 46937 12795 46995 12801
rect 47029 12835 47087 12841
rect 47029 12801 47041 12835
rect 47075 12832 47087 12835
rect 47210 12832 47216 12844
rect 47075 12804 47216 12832
rect 47075 12801 47087 12804
rect 47029 12795 47087 12801
rect 47210 12792 47216 12804
rect 47268 12792 47274 12844
rect 48038 12832 48044 12844
rect 47999 12804 48044 12832
rect 48038 12792 48044 12804
rect 48096 12792 48102 12844
rect 48314 12792 48320 12844
rect 48372 12832 48378 12844
rect 49160 12841 49188 12872
rect 49329 12869 49341 12903
rect 49375 12900 49387 12903
rect 49786 12900 49792 12912
rect 49375 12872 49792 12900
rect 49375 12869 49387 12872
rect 49329 12863 49387 12869
rect 49786 12860 49792 12872
rect 49844 12860 49850 12912
rect 51046 12900 51074 12940
rect 53834 12928 53840 12940
rect 53892 12928 53898 12980
rect 50448 12872 51074 12900
rect 51353 12903 51411 12909
rect 48961 12835 49019 12841
rect 48961 12832 48973 12835
rect 48372 12804 48973 12832
rect 48372 12792 48378 12804
rect 48961 12801 48973 12804
rect 49007 12801 49019 12835
rect 48961 12795 49019 12801
rect 49109 12835 49188 12841
rect 49109 12801 49121 12835
rect 49155 12804 49188 12835
rect 49237 12835 49295 12841
rect 49237 12806 49249 12835
rect 49283 12806 49295 12835
rect 49155 12801 49167 12804
rect 49109 12795 49167 12801
rect 41966 12764 41972 12776
rect 41800 12736 41972 12764
rect 41966 12724 41972 12736
rect 42024 12764 42030 12776
rect 45186 12764 45192 12776
rect 42024 12736 45192 12764
rect 42024 12724 42030 12736
rect 45186 12724 45192 12736
rect 45244 12724 45250 12776
rect 46017 12767 46075 12773
rect 46017 12733 46029 12767
rect 46063 12764 46075 12767
rect 46658 12764 46664 12776
rect 46063 12736 46664 12764
rect 46063 12733 46075 12736
rect 46017 12727 46075 12733
rect 46658 12724 46664 12736
rect 46716 12724 46722 12776
rect 46750 12724 46756 12776
rect 46808 12764 46814 12776
rect 46808 12736 46853 12764
rect 49234 12754 49240 12806
rect 49292 12754 49298 12806
rect 49418 12792 49424 12844
rect 49476 12841 49482 12844
rect 49476 12832 49484 12841
rect 50448 12832 50476 12872
rect 51353 12869 51365 12903
rect 51399 12900 51411 12903
rect 52086 12900 52092 12912
rect 51399 12872 52092 12900
rect 51399 12869 51411 12872
rect 51353 12863 51411 12869
rect 52086 12860 52092 12872
rect 52144 12860 52150 12912
rect 52546 12860 52552 12912
rect 52604 12900 52610 12912
rect 56226 12900 56232 12912
rect 52604 12872 54708 12900
rect 52604 12860 52610 12872
rect 50614 12832 50620 12844
rect 49476 12804 50476 12832
rect 50575 12804 50620 12832
rect 49476 12795 49484 12804
rect 49476 12792 49482 12795
rect 50614 12792 50620 12804
rect 50672 12792 50678 12844
rect 50801 12835 50859 12841
rect 50801 12801 50813 12835
rect 50847 12832 50859 12835
rect 51902 12832 51908 12844
rect 50847 12804 51908 12832
rect 50847 12801 50859 12804
rect 50801 12795 50859 12801
rect 51902 12792 51908 12804
rect 51960 12792 51966 12844
rect 52181 12835 52239 12841
rect 52181 12801 52193 12835
rect 52227 12801 52239 12835
rect 52181 12795 52239 12801
rect 52365 12835 52423 12841
rect 52365 12801 52377 12835
rect 52411 12832 52423 12835
rect 52454 12832 52460 12844
rect 52411 12804 52460 12832
rect 52411 12801 52423 12804
rect 52365 12795 52423 12801
rect 49786 12764 49792 12776
rect 49344 12736 49792 12764
rect 46808 12724 46814 12736
rect 38764 12668 39068 12696
rect 39209 12699 39267 12705
rect 38197 12659 38255 12665
rect 39209 12665 39221 12699
rect 39255 12696 39267 12699
rect 40126 12696 40132 12708
rect 39255 12668 40132 12696
rect 39255 12665 39267 12668
rect 39209 12659 39267 12665
rect 40126 12656 40132 12668
rect 40184 12656 40190 12708
rect 40221 12699 40279 12705
rect 40221 12665 40233 12699
rect 40267 12696 40279 12699
rect 40402 12696 40408 12708
rect 40267 12668 40408 12696
rect 40267 12665 40279 12668
rect 40221 12659 40279 12665
rect 40402 12656 40408 12668
rect 40460 12656 40466 12708
rect 44542 12696 44548 12708
rect 44503 12668 44548 12696
rect 44542 12656 44548 12668
rect 44600 12656 44606 12708
rect 44634 12656 44640 12708
rect 44692 12696 44698 12708
rect 44910 12696 44916 12708
rect 44692 12668 44916 12696
rect 44692 12656 44698 12668
rect 44910 12656 44916 12668
rect 44968 12656 44974 12708
rect 37182 12628 37188 12640
rect 35176 12600 37188 12628
rect 37182 12588 37188 12600
rect 37240 12588 37246 12640
rect 39025 12631 39083 12637
rect 39025 12597 39037 12631
rect 39071 12628 39083 12631
rect 39298 12628 39304 12640
rect 39071 12600 39304 12628
rect 39071 12597 39083 12600
rect 39025 12591 39083 12597
rect 39298 12588 39304 12600
rect 39356 12588 39362 12640
rect 40034 12628 40040 12640
rect 39995 12600 40040 12628
rect 40034 12588 40040 12600
rect 40092 12588 40098 12640
rect 41969 12631 42027 12637
rect 41969 12597 41981 12631
rect 42015 12628 42027 12631
rect 43714 12628 43720 12640
rect 42015 12600 43720 12628
rect 42015 12597 42027 12600
rect 41969 12591 42027 12597
rect 43714 12588 43720 12600
rect 43772 12588 43778 12640
rect 46109 12631 46167 12637
rect 46109 12597 46121 12631
rect 46155 12628 46167 12631
rect 46382 12628 46388 12640
rect 46155 12600 46388 12628
rect 46155 12597 46167 12600
rect 46109 12591 46167 12597
rect 46382 12588 46388 12600
rect 46440 12588 46446 12640
rect 46658 12588 46664 12640
rect 46716 12628 46722 12640
rect 46845 12631 46903 12637
rect 46845 12628 46857 12631
rect 46716 12600 46857 12628
rect 46716 12588 46722 12600
rect 46845 12597 46857 12600
rect 46891 12597 46903 12631
rect 46845 12591 46903 12597
rect 48130 12588 48136 12640
rect 48188 12628 48194 12640
rect 49344 12628 49372 12736
rect 49786 12724 49792 12736
rect 49844 12764 49850 12776
rect 50982 12764 50988 12776
rect 49844 12736 50988 12764
rect 49844 12724 49850 12736
rect 50982 12724 50988 12736
rect 51040 12724 51046 12776
rect 51350 12724 51356 12776
rect 51408 12764 51414 12776
rect 52196 12764 52224 12795
rect 52454 12792 52460 12804
rect 52512 12792 52518 12844
rect 52914 12832 52920 12844
rect 52875 12804 52920 12832
rect 52914 12792 52920 12804
rect 52972 12792 52978 12844
rect 53098 12792 53104 12844
rect 53156 12832 53162 12844
rect 54680 12841 54708 12872
rect 54864 12872 56232 12900
rect 54864 12844 54892 12872
rect 56226 12860 56232 12872
rect 56284 12860 56290 12912
rect 56962 12860 56968 12912
rect 57020 12900 57026 12912
rect 57882 12900 57888 12912
rect 57020 12872 57888 12900
rect 57020 12860 57026 12872
rect 57882 12860 57888 12872
rect 57940 12900 57946 12912
rect 58069 12903 58127 12909
rect 58069 12900 58081 12903
rect 57940 12872 58081 12900
rect 57940 12860 57946 12872
rect 58069 12869 58081 12872
rect 58115 12869 58127 12903
rect 58069 12863 58127 12869
rect 53193 12835 53251 12841
rect 53193 12832 53205 12835
rect 53156 12804 53205 12832
rect 53156 12792 53162 12804
rect 53193 12801 53205 12804
rect 53239 12801 53251 12835
rect 53193 12795 53251 12801
rect 54665 12835 54723 12841
rect 54665 12801 54677 12835
rect 54711 12801 54723 12835
rect 54846 12832 54852 12844
rect 54807 12804 54852 12832
rect 54665 12795 54723 12801
rect 51408 12736 52224 12764
rect 52932 12764 52960 12792
rect 53742 12764 53748 12776
rect 52932 12736 53748 12764
rect 51408 12724 51414 12736
rect 53742 12724 53748 12736
rect 53800 12724 53806 12776
rect 54680 12764 54708 12795
rect 54846 12792 54852 12804
rect 54904 12792 54910 12844
rect 55030 12832 55036 12844
rect 54991 12804 55036 12832
rect 55030 12792 55036 12804
rect 55088 12792 55094 12844
rect 55493 12835 55551 12841
rect 55493 12801 55505 12835
rect 55539 12832 55551 12835
rect 55539 12804 56364 12832
rect 55539 12801 55551 12804
rect 55493 12795 55551 12801
rect 54938 12764 54944 12776
rect 54680 12736 54944 12764
rect 54938 12724 54944 12736
rect 54996 12724 55002 12776
rect 55766 12764 55772 12776
rect 55727 12736 55772 12764
rect 55766 12724 55772 12736
rect 55824 12724 55830 12776
rect 49970 12656 49976 12708
rect 50028 12696 50034 12708
rect 51074 12696 51080 12708
rect 50028 12668 51080 12696
rect 50028 12656 50034 12668
rect 51074 12656 51080 12668
rect 51132 12656 51138 12708
rect 52086 12656 52092 12708
rect 52144 12696 52150 12708
rect 53837 12699 53895 12705
rect 53837 12696 53849 12699
rect 52144 12668 53849 12696
rect 52144 12656 52150 12668
rect 53837 12665 53849 12668
rect 53883 12696 53895 12699
rect 54386 12696 54392 12708
rect 53883 12668 54392 12696
rect 53883 12665 53895 12668
rect 53837 12659 53895 12665
rect 54386 12656 54392 12668
rect 54444 12656 54450 12708
rect 49602 12628 49608 12640
rect 48188 12600 49372 12628
rect 49563 12600 49608 12628
rect 48188 12588 48194 12600
rect 49602 12588 49608 12600
rect 49660 12588 49666 12640
rect 52365 12631 52423 12637
rect 52365 12597 52377 12631
rect 52411 12628 52423 12631
rect 53009 12631 53067 12637
rect 53009 12628 53021 12631
rect 52411 12600 53021 12628
rect 52411 12597 52423 12600
rect 52365 12591 52423 12597
rect 53009 12597 53021 12600
rect 53055 12597 53067 12631
rect 53009 12591 53067 12597
rect 53377 12631 53435 12637
rect 53377 12597 53389 12631
rect 53423 12628 53435 12631
rect 53558 12628 53564 12640
rect 53423 12600 53564 12628
rect 53423 12597 53435 12600
rect 53377 12591 53435 12597
rect 53558 12588 53564 12600
rect 53616 12588 53622 12640
rect 55398 12588 55404 12640
rect 55456 12628 55462 12640
rect 55585 12631 55643 12637
rect 55585 12628 55597 12631
rect 55456 12600 55597 12628
rect 55456 12588 55462 12600
rect 55585 12597 55597 12600
rect 55631 12597 55643 12631
rect 55585 12591 55643 12597
rect 55674 12588 55680 12640
rect 55732 12628 55738 12640
rect 56336 12637 56364 12804
rect 56873 12699 56931 12705
rect 56873 12665 56885 12699
rect 56919 12696 56931 12699
rect 56962 12696 56968 12708
rect 56919 12668 56968 12696
rect 56919 12665 56931 12668
rect 56873 12659 56931 12665
rect 56962 12656 56968 12668
rect 57020 12656 57026 12708
rect 56321 12631 56379 12637
rect 55732 12600 55777 12628
rect 55732 12588 55738 12600
rect 56321 12597 56333 12631
rect 56367 12628 56379 12631
rect 56686 12628 56692 12640
rect 56367 12600 56692 12628
rect 56367 12597 56379 12600
rect 56321 12591 56379 12597
rect 56686 12588 56692 12600
rect 56744 12628 56750 12640
rect 57422 12628 57428 12640
rect 56744 12600 57428 12628
rect 56744 12588 56750 12600
rect 57422 12588 57428 12600
rect 57480 12588 57486 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 24486 12384 24492 12436
rect 24544 12424 24550 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 24544 12396 24593 12424
rect 24544 12384 24550 12396
rect 24581 12393 24593 12396
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 25774 12384 25780 12436
rect 25832 12424 25838 12436
rect 26053 12427 26111 12433
rect 26053 12424 26065 12427
rect 25832 12396 26065 12424
rect 25832 12384 25838 12396
rect 26053 12393 26065 12396
rect 26099 12393 26111 12427
rect 26053 12387 26111 12393
rect 27157 12427 27215 12433
rect 27157 12393 27169 12427
rect 27203 12424 27215 12427
rect 27430 12424 27436 12436
rect 27203 12396 27436 12424
rect 27203 12393 27215 12396
rect 27157 12387 27215 12393
rect 27430 12384 27436 12396
rect 27488 12384 27494 12436
rect 32309 12427 32367 12433
rect 27632 12396 32260 12424
rect 25501 12359 25559 12365
rect 25501 12325 25513 12359
rect 25547 12356 25559 12359
rect 25682 12356 25688 12368
rect 25547 12328 25688 12356
rect 25547 12325 25559 12328
rect 25501 12319 25559 12325
rect 25682 12316 25688 12328
rect 25740 12356 25746 12368
rect 27632 12356 27660 12396
rect 25740 12328 27660 12356
rect 25740 12316 25746 12328
rect 27338 12288 27344 12300
rect 27299 12260 27344 12288
rect 27338 12248 27344 12260
rect 27396 12248 27402 12300
rect 27430 12248 27436 12300
rect 27488 12288 27494 12300
rect 27632 12297 27660 12328
rect 28810 12316 28816 12368
rect 28868 12356 28874 12368
rect 30374 12356 30380 12368
rect 28868 12328 30380 12356
rect 28868 12316 28874 12328
rect 30374 12316 30380 12328
rect 30432 12316 30438 12368
rect 32232 12356 32260 12396
rect 32309 12393 32321 12427
rect 32355 12424 32367 12427
rect 32490 12424 32496 12436
rect 32355 12396 32496 12424
rect 32355 12393 32367 12396
rect 32309 12387 32367 12393
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 33134 12424 33140 12436
rect 33095 12396 33140 12424
rect 33134 12384 33140 12396
rect 33192 12384 33198 12436
rect 36630 12384 36636 12436
rect 36688 12424 36694 12436
rect 36725 12427 36783 12433
rect 36725 12424 36737 12427
rect 36688 12396 36737 12424
rect 36688 12384 36694 12396
rect 36725 12393 36737 12396
rect 36771 12393 36783 12427
rect 36725 12387 36783 12393
rect 37182 12384 37188 12436
rect 37240 12424 37246 12436
rect 37461 12427 37519 12433
rect 37461 12424 37473 12427
rect 37240 12396 37473 12424
rect 37240 12384 37246 12396
rect 37461 12393 37473 12396
rect 37507 12393 37519 12427
rect 38838 12424 38844 12436
rect 37461 12387 37519 12393
rect 37844 12396 38844 12424
rect 32398 12356 32404 12368
rect 32232 12328 32404 12356
rect 32398 12316 32404 12328
rect 32456 12316 32462 12368
rect 33612 12328 36308 12356
rect 27617 12291 27675 12297
rect 27488 12260 27533 12288
rect 27488 12248 27494 12260
rect 27617 12257 27629 12291
rect 27663 12257 27675 12291
rect 28828 12288 28856 12316
rect 30561 12291 30619 12297
rect 30561 12288 30573 12291
rect 27617 12251 27675 12257
rect 28552 12260 28856 12288
rect 28920 12260 30573 12288
rect 27522 12220 27528 12232
rect 27483 12192 27528 12220
rect 27522 12180 27528 12192
rect 27580 12180 27586 12232
rect 28552 12229 28580 12260
rect 28537 12223 28595 12229
rect 28537 12189 28549 12223
rect 28583 12189 28595 12223
rect 28718 12220 28724 12232
rect 28679 12192 28724 12220
rect 28537 12183 28595 12189
rect 28718 12180 28724 12192
rect 28776 12180 28782 12232
rect 28920 12229 28948 12260
rect 30561 12257 30573 12260
rect 30607 12257 30619 12291
rect 33318 12288 33324 12300
rect 33279 12260 33324 12288
rect 30561 12251 30619 12257
rect 33318 12248 33324 12260
rect 33376 12248 33382 12300
rect 28813 12223 28871 12229
rect 28813 12189 28825 12223
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 28905 12223 28963 12229
rect 28905 12189 28917 12223
rect 28951 12189 28963 12223
rect 28905 12183 28963 12189
rect 28997 12223 29055 12229
rect 28997 12189 29009 12223
rect 29043 12220 29055 12223
rect 30190 12220 30196 12232
rect 29043 12192 30196 12220
rect 29043 12189 29055 12192
rect 28997 12183 29055 12189
rect 25225 12155 25283 12161
rect 25225 12121 25237 12155
rect 25271 12152 25283 12155
rect 25271 12124 25305 12152
rect 25271 12121 25283 12124
rect 25225 12115 25283 12121
rect 24029 12087 24087 12093
rect 24029 12053 24041 12087
rect 24075 12084 24087 12087
rect 25240 12084 25268 12115
rect 26786 12112 26792 12164
rect 26844 12152 26850 12164
rect 28074 12152 28080 12164
rect 26844 12124 28080 12152
rect 26844 12112 26850 12124
rect 28074 12112 28080 12124
rect 28132 12112 28138 12164
rect 28350 12112 28356 12164
rect 28408 12152 28414 12164
rect 28828 12152 28856 12183
rect 28408 12124 28856 12152
rect 28408 12112 28414 12124
rect 26602 12084 26608 12096
rect 24075 12056 26608 12084
rect 24075 12053 24087 12056
rect 24029 12047 24087 12053
rect 26602 12044 26608 12056
rect 26660 12084 26666 12096
rect 26878 12084 26884 12096
rect 26660 12056 26884 12084
rect 26660 12044 26666 12056
rect 26878 12044 26884 12056
rect 26936 12044 26942 12096
rect 28626 12044 28632 12096
rect 28684 12084 28690 12096
rect 28920 12084 28948 12183
rect 30190 12180 30196 12192
rect 30248 12180 30254 12232
rect 30282 12180 30288 12232
rect 30340 12220 30346 12232
rect 30469 12223 30527 12229
rect 30340 12192 30385 12220
rect 30340 12180 30346 12192
rect 30469 12189 30481 12223
rect 30515 12189 30527 12223
rect 30469 12183 30527 12189
rect 30653 12223 30711 12229
rect 30653 12189 30665 12223
rect 30699 12189 30711 12223
rect 30653 12183 30711 12189
rect 30006 12112 30012 12164
rect 30064 12152 30070 12164
rect 30101 12155 30159 12161
rect 30101 12152 30113 12155
rect 30064 12124 30113 12152
rect 30064 12112 30070 12124
rect 30101 12121 30113 12124
rect 30147 12121 30159 12155
rect 30101 12115 30159 12121
rect 30374 12112 30380 12164
rect 30432 12152 30438 12164
rect 30484 12152 30512 12183
rect 30432 12124 30512 12152
rect 30668 12152 30696 12183
rect 30742 12180 30748 12232
rect 30800 12220 30806 12232
rect 30837 12223 30895 12229
rect 30837 12220 30849 12223
rect 30800 12192 30849 12220
rect 30800 12180 30806 12192
rect 30837 12189 30849 12192
rect 30883 12189 30895 12223
rect 30837 12183 30895 12189
rect 31941 12223 31999 12229
rect 31941 12189 31953 12223
rect 31987 12220 31999 12223
rect 33042 12220 33048 12232
rect 31987 12192 33048 12220
rect 31987 12189 31999 12192
rect 31941 12183 31999 12189
rect 33042 12180 33048 12192
rect 33100 12180 33106 12232
rect 33410 12180 33416 12232
rect 33468 12220 33474 12232
rect 33468 12192 33513 12220
rect 33468 12180 33474 12192
rect 31846 12152 31852 12164
rect 30668 12124 31852 12152
rect 30432 12112 30438 12124
rect 31846 12112 31852 12124
rect 31904 12112 31910 12164
rect 32125 12155 32183 12161
rect 32125 12121 32137 12155
rect 32171 12152 32183 12155
rect 33612 12152 33640 12328
rect 34422 12248 34428 12300
rect 34480 12288 34486 12300
rect 36280 12288 36308 12328
rect 37734 12288 37740 12300
rect 34480 12260 35848 12288
rect 34480 12248 34486 12260
rect 33686 12180 33692 12232
rect 33744 12220 33750 12232
rect 33744 12192 33789 12220
rect 33744 12180 33750 12192
rect 33870 12180 33876 12232
rect 33928 12220 33934 12232
rect 34885 12223 34943 12229
rect 34885 12220 34897 12223
rect 33928 12192 34897 12220
rect 33928 12180 33934 12192
rect 34885 12189 34897 12192
rect 34931 12189 34943 12223
rect 34885 12183 34943 12189
rect 35066 12180 35072 12232
rect 35124 12220 35130 12232
rect 35820 12229 35848 12260
rect 36280 12260 37740 12288
rect 36280 12229 36308 12260
rect 37734 12248 37740 12260
rect 37792 12248 37798 12300
rect 37844 12297 37872 12396
rect 38838 12384 38844 12396
rect 38896 12384 38902 12436
rect 39301 12427 39359 12433
rect 39301 12393 39313 12427
rect 39347 12424 39359 12427
rect 39390 12424 39396 12436
rect 39347 12396 39396 12424
rect 39347 12393 39359 12396
rect 39301 12387 39359 12393
rect 39390 12384 39396 12396
rect 39448 12424 39454 12436
rect 40586 12424 40592 12436
rect 39448 12396 40448 12424
rect 40547 12396 40592 12424
rect 39448 12384 39454 12396
rect 37918 12316 37924 12368
rect 37976 12356 37982 12368
rect 37976 12328 38240 12356
rect 37976 12316 37982 12328
rect 37829 12291 37887 12297
rect 37829 12257 37841 12291
rect 37875 12257 37887 12291
rect 37829 12251 37887 12257
rect 35621 12223 35679 12229
rect 35621 12220 35633 12223
rect 35124 12192 35633 12220
rect 35124 12180 35130 12192
rect 35621 12189 35633 12192
rect 35667 12189 35679 12223
rect 35621 12183 35679 12189
rect 35805 12223 35863 12229
rect 35805 12189 35817 12223
rect 35851 12189 35863 12223
rect 35805 12183 35863 12189
rect 36265 12223 36323 12229
rect 36265 12189 36277 12223
rect 36311 12189 36323 12223
rect 36265 12183 36323 12189
rect 36354 12180 36360 12232
rect 36412 12220 36418 12232
rect 36541 12223 36599 12229
rect 36541 12220 36553 12223
rect 36412 12192 36553 12220
rect 36412 12180 36418 12192
rect 36541 12189 36553 12192
rect 36587 12220 36599 12223
rect 36722 12220 36728 12232
rect 36587 12192 36728 12220
rect 36587 12189 36599 12192
rect 36541 12183 36599 12189
rect 36722 12180 36728 12192
rect 36780 12220 36786 12232
rect 37642 12220 37648 12232
rect 36780 12192 37412 12220
rect 37603 12192 37648 12220
rect 36780 12180 36786 12192
rect 32171 12124 33640 12152
rect 32171 12121 32183 12124
rect 32125 12115 32183 12121
rect 28684 12056 28948 12084
rect 29181 12087 29239 12093
rect 28684 12044 28690 12056
rect 29181 12053 29193 12087
rect 29227 12084 29239 12087
rect 29270 12084 29276 12096
rect 29227 12056 29276 12084
rect 29227 12053 29239 12056
rect 29181 12047 29239 12053
rect 29270 12044 29276 12056
rect 29328 12044 29334 12096
rect 30742 12044 30748 12096
rect 30800 12084 30806 12096
rect 31938 12084 31944 12096
rect 30800 12056 31944 12084
rect 30800 12044 30806 12056
rect 31938 12044 31944 12056
rect 31996 12084 32002 12096
rect 32140 12084 32168 12115
rect 33778 12112 33784 12164
rect 33836 12152 33842 12164
rect 33836 12124 33881 12152
rect 33836 12112 33842 12124
rect 34054 12112 34060 12164
rect 34112 12152 34118 12164
rect 34977 12155 35035 12161
rect 34977 12152 34989 12155
rect 34112 12124 34989 12152
rect 34112 12112 34118 12124
rect 34977 12121 34989 12124
rect 35023 12121 35035 12155
rect 34977 12115 35035 12121
rect 35161 12155 35219 12161
rect 35161 12121 35173 12155
rect 35207 12152 35219 12155
rect 37274 12152 37280 12164
rect 35207 12124 37280 12152
rect 35207 12121 35219 12124
rect 35161 12115 35219 12121
rect 37274 12112 37280 12124
rect 37332 12112 37338 12164
rect 37384 12152 37412 12192
rect 37642 12180 37648 12192
rect 37700 12180 37706 12232
rect 37918 12220 37924 12232
rect 37879 12192 37924 12220
rect 37918 12180 37924 12192
rect 37976 12180 37982 12232
rect 38013 12223 38071 12229
rect 38013 12189 38025 12223
rect 38059 12220 38071 12223
rect 38102 12220 38108 12232
rect 38059 12192 38108 12220
rect 38059 12189 38071 12192
rect 38013 12183 38071 12189
rect 38102 12180 38108 12192
rect 38160 12180 38166 12232
rect 38212 12229 38240 12328
rect 40034 12316 40040 12368
rect 40092 12356 40098 12368
rect 40221 12359 40279 12365
rect 40221 12356 40233 12359
rect 40092 12328 40233 12356
rect 40092 12316 40098 12328
rect 40221 12325 40233 12328
rect 40267 12325 40279 12359
rect 40420 12356 40448 12396
rect 40586 12384 40592 12396
rect 40644 12384 40650 12436
rect 42153 12427 42211 12433
rect 42153 12424 42165 12427
rect 40696 12396 42165 12424
rect 40696 12368 40724 12396
rect 42153 12393 42165 12396
rect 42199 12393 42211 12427
rect 42153 12387 42211 12393
rect 43625 12427 43683 12433
rect 43625 12393 43637 12427
rect 43671 12424 43683 12427
rect 44082 12424 44088 12436
rect 43671 12396 44088 12424
rect 43671 12393 43683 12396
rect 43625 12387 43683 12393
rect 44082 12384 44088 12396
rect 44140 12384 44146 12436
rect 46106 12384 46112 12436
rect 46164 12424 46170 12436
rect 46385 12427 46443 12433
rect 46385 12424 46397 12427
rect 46164 12396 46397 12424
rect 46164 12384 46170 12396
rect 46385 12393 46397 12396
rect 46431 12393 46443 12427
rect 46385 12387 46443 12393
rect 48130 12384 48136 12436
rect 48188 12424 48194 12436
rect 48590 12424 48596 12436
rect 48188 12396 48596 12424
rect 48188 12384 48194 12396
rect 48590 12384 48596 12396
rect 48648 12384 48654 12436
rect 48774 12384 48780 12436
rect 48832 12424 48838 12436
rect 49513 12427 49571 12433
rect 49513 12424 49525 12427
rect 48832 12396 49525 12424
rect 48832 12384 48838 12396
rect 49513 12393 49525 12396
rect 49559 12393 49571 12427
rect 49513 12387 49571 12393
rect 50706 12384 50712 12436
rect 50764 12424 50770 12436
rect 52086 12424 52092 12436
rect 50764 12396 52092 12424
rect 50764 12384 50770 12396
rect 52086 12384 52092 12396
rect 52144 12384 52150 12436
rect 52917 12427 52975 12433
rect 52917 12393 52929 12427
rect 52963 12424 52975 12427
rect 53561 12427 53619 12433
rect 53561 12424 53573 12427
rect 52963 12396 53573 12424
rect 52963 12393 52975 12396
rect 52917 12387 52975 12393
rect 53561 12393 53573 12396
rect 53607 12393 53619 12427
rect 53561 12387 53619 12393
rect 53650 12384 53656 12436
rect 53708 12384 53714 12436
rect 54018 12384 54024 12436
rect 54076 12424 54082 12436
rect 54389 12427 54447 12433
rect 54389 12424 54401 12427
rect 54076 12396 54401 12424
rect 54076 12384 54082 12396
rect 54389 12393 54401 12396
rect 54435 12393 54447 12427
rect 54389 12387 54447 12393
rect 54938 12384 54944 12436
rect 54996 12424 55002 12436
rect 56689 12427 56747 12433
rect 56689 12424 56701 12427
rect 54996 12396 56701 12424
rect 54996 12384 55002 12396
rect 56689 12393 56701 12396
rect 56735 12424 56747 12427
rect 58066 12424 58072 12436
rect 56735 12396 58072 12424
rect 56735 12393 56747 12396
rect 56689 12387 56747 12393
rect 58066 12384 58072 12396
rect 58124 12384 58130 12436
rect 40678 12356 40684 12368
rect 40420 12328 40684 12356
rect 40221 12319 40279 12325
rect 40678 12316 40684 12328
rect 40736 12316 40742 12368
rect 43162 12316 43168 12368
rect 43220 12356 43226 12368
rect 43714 12356 43720 12368
rect 43220 12328 43720 12356
rect 43220 12316 43226 12328
rect 43714 12316 43720 12328
rect 43772 12316 43778 12368
rect 44910 12316 44916 12368
rect 44968 12356 44974 12368
rect 45189 12359 45247 12365
rect 45189 12356 45201 12359
rect 44968 12328 45201 12356
rect 44968 12316 44974 12328
rect 45189 12325 45201 12328
rect 45235 12325 45247 12359
rect 45189 12319 45247 12325
rect 45278 12316 45284 12368
rect 45336 12356 45342 12368
rect 47489 12359 47547 12365
rect 47489 12356 47501 12359
rect 45336 12328 47501 12356
rect 45336 12316 45342 12328
rect 47489 12325 47501 12328
rect 47535 12356 47547 12359
rect 48314 12356 48320 12368
rect 47535 12328 48320 12356
rect 47535 12325 47547 12328
rect 47489 12319 47547 12325
rect 48314 12316 48320 12328
rect 48372 12316 48378 12368
rect 48498 12356 48504 12368
rect 48424 12328 48504 12356
rect 43530 12288 43536 12300
rect 42996 12260 43536 12288
rect 38197 12223 38255 12229
rect 38197 12189 38209 12223
rect 38243 12189 38255 12223
rect 40126 12220 40132 12232
rect 40087 12192 40132 12220
rect 38197 12183 38255 12189
rect 40126 12180 40132 12192
rect 40184 12180 40190 12232
rect 40310 12220 40316 12232
rect 40271 12192 40316 12220
rect 40310 12180 40316 12192
rect 40368 12180 40374 12232
rect 40402 12180 40408 12232
rect 40460 12220 40466 12232
rect 42996 12229 43024 12260
rect 43530 12248 43536 12260
rect 43588 12248 43594 12300
rect 45554 12248 45560 12300
rect 45612 12288 45618 12300
rect 45922 12288 45928 12300
rect 45612 12260 45928 12288
rect 45612 12248 45618 12260
rect 45922 12248 45928 12260
rect 45980 12248 45986 12300
rect 48130 12288 48136 12300
rect 46768 12260 48136 12288
rect 42981 12223 43039 12229
rect 40460 12192 40505 12220
rect 40460 12180 40466 12192
rect 42981 12189 42993 12223
rect 43027 12189 43039 12223
rect 43162 12220 43168 12232
rect 43123 12192 43168 12220
rect 42981 12183 43039 12189
rect 38657 12155 38715 12161
rect 38657 12152 38669 12155
rect 37384 12124 38669 12152
rect 38657 12121 38669 12124
rect 38703 12121 38715 12155
rect 42996 12152 43024 12183
rect 43162 12180 43168 12192
rect 43220 12180 43226 12232
rect 43260 12223 43318 12229
rect 43260 12220 43272 12223
rect 43259 12189 43272 12220
rect 43306 12189 43318 12223
rect 43259 12183 43318 12189
rect 43070 12152 43076 12164
rect 42996 12124 43076 12152
rect 38657 12115 38715 12121
rect 43070 12112 43076 12124
rect 43128 12112 43134 12164
rect 43259 12096 43287 12183
rect 43346 12180 43352 12232
rect 43404 12220 43410 12232
rect 43404 12192 43449 12220
rect 43404 12180 43410 12192
rect 45462 12180 45468 12232
rect 45520 12220 45526 12232
rect 46768 12229 46796 12260
rect 48130 12248 48136 12260
rect 48188 12248 48194 12300
rect 48424 12288 48452 12328
rect 48498 12316 48504 12328
rect 48556 12316 48562 12368
rect 49418 12316 49424 12368
rect 49476 12356 49482 12368
rect 52641 12359 52699 12365
rect 49476 12328 51580 12356
rect 49476 12316 49482 12328
rect 48958 12288 48964 12300
rect 48332 12260 48452 12288
rect 48516 12260 48964 12288
rect 46569 12223 46627 12229
rect 46569 12220 46581 12223
rect 45520 12192 45565 12220
rect 46492 12192 46581 12220
rect 45520 12180 45526 12192
rect 43990 12112 43996 12164
rect 44048 12152 44054 12164
rect 45189 12155 45247 12161
rect 45189 12152 45201 12155
rect 44048 12124 45201 12152
rect 44048 12112 44054 12124
rect 45189 12121 45201 12124
rect 45235 12121 45247 12155
rect 45189 12115 45247 12121
rect 45278 12112 45284 12164
rect 45336 12152 45342 12164
rect 45646 12152 45652 12164
rect 45336 12124 45652 12152
rect 45336 12112 45342 12124
rect 45646 12112 45652 12124
rect 45704 12112 45710 12164
rect 46106 12112 46112 12164
rect 46164 12152 46170 12164
rect 46290 12152 46296 12164
rect 46164 12124 46296 12152
rect 46164 12112 46170 12124
rect 46290 12112 46296 12124
rect 46348 12112 46354 12164
rect 31996 12056 32168 12084
rect 31996 12044 32002 12056
rect 32398 12044 32404 12096
rect 32456 12084 32462 12096
rect 34241 12087 34299 12093
rect 34241 12084 34253 12087
rect 32456 12056 34253 12084
rect 32456 12044 32462 12056
rect 34241 12053 34253 12056
rect 34287 12084 34299 12087
rect 34882 12084 34888 12096
rect 34287 12056 34888 12084
rect 34287 12053 34299 12056
rect 34241 12047 34299 12053
rect 34882 12044 34888 12056
rect 34940 12044 34946 12096
rect 35062 12087 35120 12093
rect 35062 12053 35074 12087
rect 35108 12084 35120 12087
rect 35250 12084 35256 12096
rect 35108 12056 35256 12084
rect 35108 12053 35120 12056
rect 35062 12047 35120 12053
rect 35250 12044 35256 12056
rect 35308 12044 35314 12096
rect 35713 12087 35771 12093
rect 35713 12053 35725 12087
rect 35759 12084 35771 12087
rect 35894 12084 35900 12096
rect 35759 12056 35900 12084
rect 35759 12053 35771 12056
rect 35713 12047 35771 12053
rect 35894 12044 35900 12056
rect 35952 12084 35958 12096
rect 36170 12084 36176 12096
rect 35952 12056 36176 12084
rect 35952 12044 35958 12056
rect 36170 12044 36176 12056
rect 36228 12044 36234 12096
rect 36357 12087 36415 12093
rect 36357 12053 36369 12087
rect 36403 12084 36415 12087
rect 36630 12084 36636 12096
rect 36403 12056 36636 12084
rect 36403 12053 36415 12056
rect 36357 12047 36415 12053
rect 36630 12044 36636 12056
rect 36688 12084 36694 12096
rect 36814 12084 36820 12096
rect 36688 12056 36820 12084
rect 36688 12044 36694 12056
rect 36814 12044 36820 12056
rect 36872 12084 36878 12096
rect 37642 12084 37648 12096
rect 36872 12056 37648 12084
rect 36872 12044 36878 12056
rect 37642 12044 37648 12056
rect 37700 12044 37706 12096
rect 38102 12044 38108 12096
rect 38160 12084 38166 12096
rect 38562 12084 38568 12096
rect 38160 12056 38568 12084
rect 38160 12044 38166 12056
rect 38562 12044 38568 12056
rect 38620 12044 38626 12096
rect 40954 12044 40960 12096
rect 41012 12084 41018 12096
rect 41049 12087 41107 12093
rect 41049 12084 41061 12087
rect 41012 12056 41061 12084
rect 41012 12044 41018 12056
rect 41049 12053 41061 12056
rect 41095 12053 41107 12087
rect 41049 12047 41107 12053
rect 41230 12044 41236 12096
rect 41288 12084 41294 12096
rect 41601 12087 41659 12093
rect 41601 12084 41613 12087
rect 41288 12056 41613 12084
rect 41288 12044 41294 12056
rect 41601 12053 41613 12056
rect 41647 12053 41659 12087
rect 41601 12047 41659 12053
rect 43254 12044 43260 12096
rect 43312 12044 43318 12096
rect 44174 12084 44180 12096
rect 44135 12056 44180 12084
rect 44174 12044 44180 12056
rect 44232 12044 44238 12096
rect 45373 12087 45431 12093
rect 45373 12053 45385 12087
rect 45419 12084 45431 12087
rect 45462 12084 45468 12096
rect 45419 12056 45468 12084
rect 45419 12053 45431 12056
rect 45373 12047 45431 12053
rect 45462 12044 45468 12056
rect 45520 12044 45526 12096
rect 45554 12044 45560 12096
rect 45612 12084 45618 12096
rect 46492 12084 46520 12192
rect 46569 12189 46581 12192
rect 46615 12189 46627 12223
rect 46569 12183 46627 12189
rect 46753 12223 46811 12229
rect 46753 12189 46765 12223
rect 46799 12189 46811 12223
rect 47026 12220 47032 12232
rect 46987 12192 47032 12220
rect 46753 12183 46811 12189
rect 47026 12180 47032 12192
rect 47084 12180 47090 12232
rect 48225 12223 48283 12229
rect 48225 12189 48237 12223
rect 48271 12189 48283 12223
rect 48332 12220 48360 12260
rect 48516 12229 48544 12260
rect 48958 12248 48964 12260
rect 49016 12248 49022 12300
rect 49694 12288 49700 12300
rect 49436 12260 49700 12288
rect 48388 12223 48446 12229
rect 48388 12220 48400 12223
rect 48332 12192 48400 12220
rect 48225 12183 48283 12189
rect 48388 12189 48400 12192
rect 48434 12189 48446 12223
rect 48388 12183 48446 12189
rect 48488 12223 48546 12229
rect 48488 12189 48500 12223
rect 48534 12189 48546 12223
rect 48488 12183 48546 12189
rect 46658 12152 46664 12164
rect 46619 12124 46664 12152
rect 46658 12112 46664 12124
rect 46716 12112 46722 12164
rect 46842 12112 46848 12164
rect 46900 12161 46906 12164
rect 46900 12155 46929 12161
rect 46917 12121 46929 12155
rect 46900 12115 46929 12121
rect 46900 12112 46906 12115
rect 47118 12112 47124 12164
rect 47176 12152 47182 12164
rect 48240 12152 48268 12183
rect 48590 12180 48596 12232
rect 48648 12220 48654 12232
rect 49436 12229 49464 12260
rect 49694 12248 49700 12260
rect 49752 12248 49758 12300
rect 50338 12248 50344 12300
rect 50396 12288 50402 12300
rect 50709 12291 50767 12297
rect 50709 12288 50721 12291
rect 50396 12260 50721 12288
rect 50396 12248 50402 12260
rect 50709 12257 50721 12260
rect 50755 12257 50767 12291
rect 50709 12251 50767 12257
rect 50801 12291 50859 12297
rect 50801 12257 50813 12291
rect 50847 12288 50859 12291
rect 50908 12288 50936 12328
rect 51552 12297 51580 12328
rect 52641 12325 52653 12359
rect 52687 12356 52699 12359
rect 52730 12356 52736 12368
rect 52687 12328 52736 12356
rect 52687 12325 52699 12328
rect 52641 12319 52699 12325
rect 52730 12316 52736 12328
rect 52788 12316 52794 12368
rect 53374 12356 53380 12368
rect 53335 12328 53380 12356
rect 53374 12316 53380 12328
rect 53432 12316 53438 12368
rect 53668 12356 53696 12384
rect 54478 12356 54484 12368
rect 53668 12328 54484 12356
rect 54478 12316 54484 12328
rect 54536 12316 54542 12368
rect 55490 12356 55496 12368
rect 55451 12328 55496 12356
rect 55490 12316 55496 12328
rect 55548 12316 55554 12368
rect 50847 12260 50936 12288
rect 51537 12291 51595 12297
rect 50847 12257 50859 12260
rect 50801 12251 50859 12257
rect 51537 12257 51549 12291
rect 51583 12288 51595 12291
rect 51583 12260 52684 12288
rect 51583 12257 51595 12260
rect 51537 12251 51595 12257
rect 49421 12223 49479 12229
rect 48648 12192 49372 12220
rect 48648 12180 48654 12192
rect 48958 12152 48964 12164
rect 47176 12124 48964 12152
rect 47176 12112 47182 12124
rect 48958 12112 48964 12124
rect 49016 12112 49022 12164
rect 49344 12152 49372 12192
rect 49421 12189 49433 12223
rect 49467 12189 49479 12223
rect 49602 12220 49608 12232
rect 49563 12192 49608 12220
rect 49421 12183 49479 12189
rect 49602 12180 49608 12192
rect 49660 12180 49666 12232
rect 49970 12180 49976 12232
rect 50028 12220 50034 12232
rect 50525 12223 50583 12229
rect 50525 12220 50537 12223
rect 50028 12192 50537 12220
rect 50028 12180 50034 12192
rect 50525 12189 50537 12192
rect 50571 12189 50583 12223
rect 50893 12223 50951 12229
rect 50893 12220 50905 12223
rect 50525 12183 50583 12189
rect 50632 12192 50905 12220
rect 50430 12152 50436 12164
rect 49344 12124 50436 12152
rect 50430 12112 50436 12124
rect 50488 12152 50494 12164
rect 50632 12152 50660 12192
rect 50893 12189 50905 12192
rect 50939 12189 50951 12223
rect 50893 12183 50951 12189
rect 51077 12223 51135 12229
rect 51077 12189 51089 12223
rect 51123 12220 51135 12223
rect 52178 12220 52184 12232
rect 51123 12192 52184 12220
rect 51123 12189 51135 12192
rect 51077 12183 51135 12189
rect 52178 12180 52184 12192
rect 52236 12180 52242 12232
rect 52273 12223 52331 12229
rect 52273 12189 52285 12223
rect 52319 12189 52331 12223
rect 52273 12183 52331 12189
rect 50488 12124 50660 12152
rect 50488 12112 50494 12124
rect 51626 12112 51632 12164
rect 51684 12152 51690 12164
rect 52288 12152 52316 12183
rect 52362 12180 52368 12232
rect 52420 12218 52426 12232
rect 52457 12223 52515 12229
rect 52457 12218 52469 12223
rect 52420 12190 52469 12218
rect 52420 12180 52426 12190
rect 52457 12189 52469 12190
rect 52503 12189 52515 12223
rect 52457 12183 52515 12189
rect 52546 12180 52552 12232
rect 52604 12220 52610 12232
rect 52656 12220 52684 12260
rect 53282 12248 53288 12300
rect 53340 12288 53346 12300
rect 53650 12288 53656 12300
rect 53340 12260 53656 12288
rect 53340 12248 53346 12260
rect 53650 12248 53656 12260
rect 53708 12248 53714 12300
rect 55950 12248 55956 12300
rect 56008 12288 56014 12300
rect 56045 12291 56103 12297
rect 56045 12288 56057 12291
rect 56008 12260 56057 12288
rect 56008 12248 56014 12260
rect 56045 12257 56057 12260
rect 56091 12257 56103 12291
rect 56045 12251 56103 12257
rect 52733 12223 52791 12229
rect 52604 12192 52697 12220
rect 52604 12190 52684 12192
rect 52604 12180 52610 12190
rect 52733 12189 52745 12223
rect 52779 12220 52791 12223
rect 52822 12220 52828 12232
rect 52779 12192 52828 12220
rect 52779 12189 52791 12192
rect 52733 12183 52791 12189
rect 52822 12180 52828 12192
rect 52880 12180 52886 12232
rect 53558 12220 53564 12232
rect 53519 12192 53564 12220
rect 53558 12180 53564 12192
rect 53616 12180 53622 12232
rect 53834 12180 53840 12232
rect 53892 12220 53898 12232
rect 53929 12223 53987 12229
rect 53929 12220 53941 12223
rect 53892 12192 53941 12220
rect 53892 12180 53898 12192
rect 53929 12189 53941 12192
rect 53975 12189 53987 12223
rect 53929 12183 53987 12189
rect 54573 12223 54631 12229
rect 54573 12189 54585 12223
rect 54619 12220 54631 12223
rect 54662 12220 54668 12232
rect 54619 12192 54668 12220
rect 54619 12189 54631 12192
rect 54573 12183 54631 12189
rect 54662 12180 54668 12192
rect 54720 12180 54726 12232
rect 54849 12223 54907 12229
rect 54849 12189 54861 12223
rect 54895 12220 54907 12223
rect 55214 12220 55220 12232
rect 54895 12192 55220 12220
rect 54895 12189 54907 12192
rect 54849 12183 54907 12189
rect 52914 12152 52920 12164
rect 51684 12124 52920 12152
rect 51684 12112 51690 12124
rect 52914 12112 52920 12124
rect 52972 12112 52978 12164
rect 54864 12152 54892 12183
rect 55214 12180 55220 12192
rect 55272 12180 55278 12232
rect 55674 12180 55680 12232
rect 55732 12220 55738 12232
rect 55861 12223 55919 12229
rect 55861 12220 55873 12223
rect 55732 12192 55873 12220
rect 55732 12180 55738 12192
rect 55861 12189 55873 12192
rect 55907 12189 55919 12223
rect 55861 12183 55919 12189
rect 53576 12124 54892 12152
rect 53576 12096 53604 12124
rect 55490 12112 55496 12164
rect 55548 12152 55554 12164
rect 57793 12155 57851 12161
rect 57793 12152 57805 12155
rect 55548 12124 57805 12152
rect 55548 12112 55554 12124
rect 57793 12121 57805 12124
rect 57839 12121 57851 12155
rect 57793 12115 57851 12121
rect 45612 12056 46520 12084
rect 45612 12044 45618 12056
rect 48222 12044 48228 12096
rect 48280 12084 48286 12096
rect 48590 12084 48596 12096
rect 48280 12056 48596 12084
rect 48280 12044 48286 12056
rect 48590 12044 48596 12056
rect 48648 12044 48654 12096
rect 48869 12087 48927 12093
rect 48869 12053 48881 12087
rect 48915 12084 48927 12087
rect 49418 12084 49424 12096
rect 48915 12056 49424 12084
rect 48915 12053 48927 12056
rect 48869 12047 48927 12053
rect 49418 12044 49424 12056
rect 49476 12044 49482 12096
rect 50341 12087 50399 12093
rect 50341 12053 50353 12087
rect 50387 12084 50399 12087
rect 50798 12084 50804 12096
rect 50387 12056 50804 12084
rect 50387 12053 50399 12056
rect 50341 12047 50399 12053
rect 50798 12044 50804 12056
rect 50856 12044 50862 12096
rect 53558 12044 53564 12096
rect 53616 12044 53622 12096
rect 54202 12044 54208 12096
rect 54260 12084 54266 12096
rect 54757 12087 54815 12093
rect 54757 12084 54769 12087
rect 54260 12056 54769 12084
rect 54260 12044 54266 12056
rect 54757 12053 54769 12056
rect 54803 12084 54815 12087
rect 54846 12084 54852 12096
rect 54803 12056 54852 12084
rect 54803 12053 54815 12056
rect 54757 12047 54815 12053
rect 54846 12044 54852 12056
rect 54904 12084 54910 12096
rect 55306 12084 55312 12096
rect 54904 12056 55312 12084
rect 54904 12044 54910 12056
rect 55306 12044 55312 12056
rect 55364 12044 55370 12096
rect 55674 12044 55680 12096
rect 55732 12084 55738 12096
rect 55953 12087 56011 12093
rect 55953 12084 55965 12087
rect 55732 12056 55965 12084
rect 55732 12044 55738 12056
rect 55953 12053 55965 12056
rect 55999 12053 56011 12087
rect 57330 12084 57336 12096
rect 57291 12056 57336 12084
rect 55953 12047 56011 12053
rect 57330 12044 57336 12056
rect 57388 12044 57394 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 24762 11880 24768 11892
rect 24723 11852 24768 11880
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 24946 11840 24952 11892
rect 25004 11880 25010 11892
rect 25501 11883 25559 11889
rect 25501 11880 25513 11883
rect 25004 11852 25513 11880
rect 25004 11840 25010 11852
rect 25501 11849 25513 11852
rect 25547 11849 25559 11883
rect 27525 11883 27583 11889
rect 27525 11880 27537 11883
rect 25501 11843 25559 11849
rect 25976 11852 27537 11880
rect 24026 11772 24032 11824
rect 24084 11812 24090 11824
rect 24121 11815 24179 11821
rect 24121 11812 24133 11815
rect 24084 11784 24133 11812
rect 24084 11772 24090 11784
rect 24121 11781 24133 11784
rect 24167 11812 24179 11815
rect 24167 11784 25176 11812
rect 24167 11781 24179 11784
rect 24121 11775 24179 11781
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 24857 11747 24915 11753
rect 1903 11716 2452 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 1670 11608 1676 11620
rect 1631 11580 1676 11608
rect 1670 11568 1676 11580
rect 1728 11568 1734 11620
rect 2424 11617 2452 11716
rect 24857 11713 24869 11747
rect 24903 11744 24915 11747
rect 24946 11744 24952 11756
rect 24903 11716 24952 11744
rect 24903 11713 24915 11716
rect 24857 11707 24915 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 25041 11747 25099 11753
rect 25041 11713 25053 11747
rect 25087 11713 25099 11747
rect 25148 11744 25176 11784
rect 25222 11772 25228 11824
rect 25280 11812 25286 11824
rect 25976 11812 26004 11852
rect 27525 11849 27537 11852
rect 27571 11880 27583 11883
rect 27890 11880 27896 11892
rect 27571 11852 27896 11880
rect 27571 11849 27583 11852
rect 27525 11843 27583 11849
rect 27890 11840 27896 11852
rect 27948 11840 27954 11892
rect 29178 11880 29184 11892
rect 29139 11852 29184 11880
rect 29178 11840 29184 11852
rect 29236 11840 29242 11892
rect 31573 11883 31631 11889
rect 31573 11849 31585 11883
rect 31619 11880 31631 11883
rect 33410 11880 33416 11892
rect 31619 11852 33416 11880
rect 31619 11849 31631 11852
rect 31573 11843 31631 11849
rect 33410 11840 33416 11852
rect 33468 11840 33474 11892
rect 33505 11883 33563 11889
rect 33505 11849 33517 11883
rect 33551 11880 33563 11883
rect 33778 11880 33784 11892
rect 33551 11852 33784 11880
rect 33551 11849 33563 11852
rect 33505 11843 33563 11849
rect 33778 11840 33784 11852
rect 33836 11840 33842 11892
rect 34054 11840 34060 11892
rect 34112 11880 34118 11892
rect 34112 11852 34192 11880
rect 34112 11840 34118 11852
rect 27154 11812 27160 11824
rect 25280 11784 26004 11812
rect 27115 11784 27160 11812
rect 25280 11772 25286 11784
rect 27154 11772 27160 11784
rect 27212 11772 27218 11824
rect 28074 11772 28080 11824
rect 28132 11812 28138 11824
rect 30837 11815 30895 11821
rect 30837 11812 30849 11815
rect 28132 11784 30849 11812
rect 28132 11772 28138 11784
rect 30837 11781 30849 11784
rect 30883 11781 30895 11815
rect 31018 11812 31024 11824
rect 30979 11784 31024 11812
rect 30837 11775 30895 11781
rect 31018 11772 31024 11784
rect 31076 11772 31082 11824
rect 31846 11772 31852 11824
rect 31904 11812 31910 11824
rect 32401 11815 32459 11821
rect 32401 11812 32413 11815
rect 31904 11784 32413 11812
rect 31904 11772 31910 11784
rect 32401 11781 32413 11784
rect 32447 11812 32459 11815
rect 33870 11812 33876 11824
rect 32447 11784 33876 11812
rect 32447 11781 32459 11784
rect 32401 11775 32459 11781
rect 33870 11772 33876 11784
rect 33928 11772 33934 11824
rect 34164 11812 34192 11852
rect 35802 11840 35808 11892
rect 35860 11880 35866 11892
rect 35860 11852 37320 11880
rect 35860 11840 35866 11852
rect 34330 11812 34336 11824
rect 34164 11784 34336 11812
rect 25682 11744 25688 11756
rect 25148 11716 25688 11744
rect 25041 11707 25099 11713
rect 2409 11611 2467 11617
rect 2409 11577 2421 11611
rect 2455 11608 2467 11611
rect 24394 11608 24400 11620
rect 2455 11580 24400 11608
rect 2455 11577 2467 11580
rect 2409 11571 2467 11577
rect 24394 11568 24400 11580
rect 24452 11568 24458 11620
rect 25056 11608 25084 11707
rect 25682 11704 25688 11716
rect 25740 11704 25746 11756
rect 26050 11744 26056 11756
rect 26011 11716 26056 11744
rect 26050 11704 26056 11716
rect 26108 11704 26114 11756
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11744 26295 11747
rect 27430 11744 27436 11756
rect 26283 11716 27436 11744
rect 26283 11713 26295 11716
rect 26237 11707 26295 11713
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 27617 11747 27675 11753
rect 27617 11713 27629 11747
rect 27663 11744 27675 11747
rect 28258 11744 28264 11756
rect 27663 11716 28264 11744
rect 27663 11713 27675 11716
rect 27617 11707 27675 11713
rect 28258 11704 28264 11716
rect 28316 11704 28322 11756
rect 28534 11704 28540 11756
rect 28592 11744 28598 11756
rect 28905 11747 28963 11753
rect 28905 11744 28917 11747
rect 28592 11716 28917 11744
rect 28592 11704 28598 11716
rect 28905 11713 28917 11716
rect 28951 11713 28963 11747
rect 29270 11744 29276 11756
rect 29231 11716 29276 11744
rect 28905 11707 28963 11713
rect 29270 11704 29276 11716
rect 29328 11704 29334 11756
rect 30742 11744 30748 11756
rect 30703 11716 30748 11744
rect 30742 11704 30748 11716
rect 30800 11704 30806 11756
rect 31481 11747 31539 11753
rect 31481 11746 31493 11747
rect 31404 11744 31493 11746
rect 30944 11718 31493 11744
rect 30944 11716 31432 11718
rect 25866 11676 25872 11688
rect 25827 11648 25872 11676
rect 25866 11636 25872 11648
rect 25924 11636 25930 11688
rect 25961 11679 26019 11685
rect 25961 11645 25973 11679
rect 26007 11676 26019 11679
rect 26418 11676 26424 11688
rect 26007 11648 26424 11676
rect 26007 11645 26019 11648
rect 25961 11639 26019 11645
rect 26418 11636 26424 11648
rect 26476 11676 26482 11688
rect 27154 11676 27160 11688
rect 26476 11648 27160 11676
rect 26476 11636 26482 11648
rect 27154 11636 27160 11648
rect 27212 11636 27218 11688
rect 27249 11679 27307 11685
rect 27249 11645 27261 11679
rect 27295 11676 27307 11679
rect 27522 11676 27528 11688
rect 27295 11648 27528 11676
rect 27295 11645 27307 11648
rect 27249 11639 27307 11645
rect 26234 11608 26240 11620
rect 25056 11580 26240 11608
rect 26234 11568 26240 11580
rect 26292 11568 26298 11620
rect 26510 11568 26516 11620
rect 26568 11608 26574 11620
rect 27264 11608 27292 11639
rect 27522 11636 27528 11648
rect 27580 11636 27586 11688
rect 28718 11676 28724 11688
rect 28679 11648 28724 11676
rect 28718 11636 28724 11648
rect 28776 11636 28782 11688
rect 30558 11636 30564 11688
rect 30616 11676 30622 11688
rect 30944 11676 30972 11716
rect 31481 11713 31493 11718
rect 31527 11713 31539 11747
rect 31481 11707 31539 11713
rect 31665 11747 31723 11753
rect 31665 11713 31677 11747
rect 31711 11713 31723 11747
rect 32490 11744 32496 11756
rect 31665 11707 31723 11713
rect 32309 11737 32367 11743
rect 30616 11648 30972 11676
rect 30616 11636 30622 11648
rect 31021 11611 31079 11617
rect 31021 11608 31033 11611
rect 26568 11580 27292 11608
rect 27356 11580 31033 11608
rect 26568 11568 26574 11580
rect 24578 11540 24584 11552
rect 24539 11512 24584 11540
rect 24578 11500 24584 11512
rect 24636 11500 24642 11552
rect 27246 11500 27252 11552
rect 27304 11540 27310 11552
rect 27356 11549 27384 11580
rect 31021 11577 31033 11580
rect 31067 11608 31079 11611
rect 31110 11608 31116 11620
rect 31067 11580 31116 11608
rect 31067 11577 31079 11580
rect 31021 11571 31079 11577
rect 31110 11568 31116 11580
rect 31168 11568 31174 11620
rect 31294 11568 31300 11620
rect 31352 11608 31358 11620
rect 31680 11608 31708 11707
rect 32309 11703 32321 11737
rect 32355 11703 32367 11737
rect 32451 11716 32496 11744
rect 32490 11704 32496 11716
rect 32548 11704 32554 11756
rect 33042 11744 33048 11756
rect 33003 11716 33048 11744
rect 33042 11704 33048 11716
rect 33100 11704 33106 11756
rect 33643 11747 33701 11753
rect 33643 11744 33655 11747
rect 33520 11716 33655 11744
rect 32309 11697 32367 11703
rect 31352 11580 31708 11608
rect 32324 11608 32352 11697
rect 33520 11688 33548 11716
rect 33643 11713 33655 11716
rect 33689 11713 33701 11747
rect 33643 11707 33701 11713
rect 33781 11747 33839 11753
rect 33781 11713 33793 11747
rect 33827 11713 33839 11747
rect 33781 11707 33839 11713
rect 33502 11636 33508 11688
rect 33560 11636 33566 11688
rect 33796 11676 33824 11707
rect 33962 11704 33968 11756
rect 34020 11744 34026 11756
rect 34164 11753 34192 11784
rect 34330 11772 34336 11784
rect 34388 11772 34394 11824
rect 35250 11812 35256 11824
rect 34716 11784 35256 11812
rect 34056 11747 34114 11753
rect 34056 11744 34068 11747
rect 34020 11716 34068 11744
rect 34020 11704 34026 11716
rect 34056 11713 34068 11716
rect 34102 11713 34114 11747
rect 34056 11707 34114 11713
rect 34149 11747 34207 11753
rect 34149 11713 34161 11747
rect 34195 11713 34207 11747
rect 34149 11707 34207 11713
rect 34238 11704 34244 11756
rect 34296 11744 34302 11756
rect 34716 11753 34744 11784
rect 35250 11772 35256 11784
rect 35308 11772 35314 11824
rect 35452 11784 36032 11812
rect 34609 11747 34667 11753
rect 34609 11744 34621 11747
rect 34296 11716 34621 11744
rect 34296 11704 34302 11716
rect 34609 11713 34621 11716
rect 34655 11713 34667 11747
rect 34609 11707 34667 11713
rect 34701 11747 34759 11753
rect 34701 11713 34713 11747
rect 34747 11713 34759 11747
rect 35452 11744 35480 11784
rect 35618 11744 35624 11756
rect 34701 11707 34759 11713
rect 34808 11716 35480 11744
rect 35579 11716 35624 11744
rect 34808 11676 34836 11716
rect 35618 11704 35624 11716
rect 35676 11704 35682 11756
rect 36004 11744 36032 11784
rect 36078 11744 36084 11756
rect 35991 11716 36084 11744
rect 36004 11714 36084 11716
rect 36078 11704 36084 11714
rect 36136 11704 36142 11756
rect 36541 11747 36599 11753
rect 36541 11713 36553 11747
rect 36587 11744 36599 11747
rect 36630 11744 36636 11756
rect 36587 11716 36636 11744
rect 36587 11713 36599 11716
rect 36541 11707 36599 11713
rect 36630 11704 36636 11716
rect 36688 11704 36694 11756
rect 36722 11704 36728 11756
rect 36780 11744 36786 11756
rect 37182 11744 37188 11756
rect 36780 11716 37188 11744
rect 36780 11704 36786 11716
rect 37182 11704 37188 11716
rect 37240 11704 37246 11756
rect 37292 11744 37320 11852
rect 37550 11840 37556 11892
rect 37608 11880 37614 11892
rect 37645 11883 37703 11889
rect 37645 11880 37657 11883
rect 37608 11852 37657 11880
rect 37608 11840 37614 11852
rect 37645 11849 37657 11852
rect 37691 11849 37703 11883
rect 37645 11843 37703 11849
rect 39393 11883 39451 11889
rect 39393 11849 39405 11883
rect 39439 11849 39451 11883
rect 39393 11843 39451 11849
rect 39022 11812 39028 11824
rect 38983 11784 39028 11812
rect 39022 11772 39028 11784
rect 39080 11772 39086 11824
rect 39114 11772 39120 11824
rect 39172 11812 39178 11824
rect 39225 11815 39283 11821
rect 39225 11812 39237 11815
rect 39172 11784 39237 11812
rect 39172 11772 39178 11784
rect 39225 11781 39237 11784
rect 39271 11781 39283 11815
rect 39408 11812 39436 11843
rect 40218 11840 40224 11892
rect 40276 11880 40282 11892
rect 40494 11880 40500 11892
rect 40276 11852 40500 11880
rect 40276 11840 40282 11852
rect 40494 11840 40500 11852
rect 40552 11880 40558 11892
rect 40681 11883 40739 11889
rect 40681 11880 40693 11883
rect 40552 11852 40693 11880
rect 40552 11840 40558 11852
rect 40681 11849 40693 11852
rect 40727 11849 40739 11883
rect 40681 11843 40739 11849
rect 42061 11883 42119 11889
rect 42061 11849 42073 11883
rect 42107 11880 42119 11883
rect 43254 11880 43260 11892
rect 42107 11852 43260 11880
rect 42107 11849 42119 11852
rect 42061 11843 42119 11849
rect 43254 11840 43260 11852
rect 43312 11840 43318 11892
rect 44266 11880 44272 11892
rect 44227 11852 44272 11880
rect 44266 11840 44272 11852
rect 44324 11840 44330 11892
rect 44453 11883 44511 11889
rect 44453 11849 44465 11883
rect 44499 11880 44511 11883
rect 45373 11883 45431 11889
rect 45373 11880 45385 11883
rect 44499 11852 45385 11880
rect 44499 11849 44511 11852
rect 44453 11843 44511 11849
rect 45373 11849 45385 11852
rect 45419 11849 45431 11883
rect 45373 11843 45431 11849
rect 45554 11840 45560 11892
rect 45612 11840 45618 11892
rect 45922 11880 45928 11892
rect 45756 11852 45928 11880
rect 40310 11812 40316 11824
rect 39408 11784 40316 11812
rect 39225 11775 39283 11781
rect 37918 11744 37924 11756
rect 37292 11716 37924 11744
rect 37918 11704 37924 11716
rect 37976 11704 37982 11756
rect 38105 11747 38163 11753
rect 38105 11713 38117 11747
rect 38151 11744 38163 11747
rect 38654 11744 38660 11756
rect 38151 11716 38660 11744
rect 38151 11713 38163 11716
rect 38105 11707 38163 11713
rect 38654 11704 38660 11716
rect 38712 11704 38718 11756
rect 40037 11747 40095 11753
rect 40037 11713 40049 11747
rect 40083 11744 40095 11747
rect 40126 11744 40132 11756
rect 40083 11716 40132 11744
rect 40083 11713 40095 11716
rect 40037 11707 40095 11713
rect 40126 11704 40132 11716
rect 40184 11704 40190 11756
rect 40236 11753 40264 11784
rect 40310 11772 40316 11784
rect 40368 11772 40374 11824
rect 43622 11812 43628 11824
rect 42352 11784 43628 11812
rect 42352 11756 42380 11784
rect 43622 11772 43628 11784
rect 43680 11772 43686 11824
rect 43717 11815 43775 11821
rect 43717 11781 43729 11815
rect 43763 11812 43775 11815
rect 45572 11812 45600 11840
rect 43763 11784 45600 11812
rect 43763 11781 43775 11784
rect 43717 11775 43775 11781
rect 40221 11747 40279 11753
rect 40221 11713 40233 11747
rect 40267 11713 40279 11747
rect 40221 11707 40279 11713
rect 41693 11747 41751 11753
rect 41693 11713 41705 11747
rect 41739 11744 41751 11747
rect 42334 11744 42340 11756
rect 41739 11716 42340 11744
rect 41739 11713 41751 11716
rect 41693 11707 41751 11713
rect 42334 11704 42340 11716
rect 42392 11704 42398 11756
rect 42978 11744 42984 11756
rect 42939 11716 42984 11744
rect 42978 11704 42984 11716
rect 43036 11704 43042 11756
rect 43070 11704 43076 11756
rect 43128 11744 43134 11756
rect 43165 11747 43223 11753
rect 43165 11744 43177 11747
rect 43128 11716 43177 11744
rect 43128 11704 43134 11716
rect 43165 11713 43177 11716
rect 43211 11713 43223 11747
rect 43438 11744 43444 11756
rect 43399 11716 43444 11744
rect 43165 11707 43223 11713
rect 43438 11704 43444 11716
rect 43496 11704 43502 11756
rect 44450 11704 44456 11756
rect 44508 11744 44514 11756
rect 44910 11744 44916 11756
rect 44508 11716 44550 11744
rect 44871 11716 44916 11744
rect 44508 11704 44514 11716
rect 44910 11704 44916 11716
rect 44968 11704 44974 11756
rect 45554 11744 45560 11756
rect 45515 11716 45560 11744
rect 45554 11704 45560 11716
rect 45612 11704 45618 11756
rect 45756 11753 45784 11852
rect 45922 11840 45928 11852
rect 45980 11880 45986 11892
rect 46290 11880 46296 11892
rect 45980 11852 46296 11880
rect 45980 11840 45986 11852
rect 46290 11840 46296 11852
rect 46348 11840 46354 11892
rect 46842 11880 46848 11892
rect 46803 11852 46848 11880
rect 46842 11840 46848 11852
rect 46900 11840 46906 11892
rect 47394 11840 47400 11892
rect 47452 11880 47458 11892
rect 47452 11852 47900 11880
rect 47452 11840 47458 11852
rect 47210 11772 47216 11824
rect 47268 11812 47274 11824
rect 47762 11812 47768 11824
rect 47268 11784 47768 11812
rect 47268 11772 47274 11784
rect 47762 11772 47768 11784
rect 47820 11772 47826 11824
rect 47872 11812 47900 11852
rect 48314 11840 48320 11892
rect 48372 11880 48378 11892
rect 48498 11880 48504 11892
rect 48372 11852 48504 11880
rect 48372 11840 48378 11852
rect 48498 11840 48504 11852
rect 48556 11840 48562 11892
rect 49142 11840 49148 11892
rect 49200 11880 49206 11892
rect 49789 11883 49847 11889
rect 49789 11880 49801 11883
rect 49200 11852 49801 11880
rect 49200 11840 49206 11852
rect 49789 11849 49801 11852
rect 49835 11849 49847 11883
rect 50614 11880 50620 11892
rect 50575 11852 50620 11880
rect 49789 11843 49847 11849
rect 50614 11840 50620 11852
rect 50672 11840 50678 11892
rect 50798 11880 50804 11892
rect 50759 11852 50804 11880
rect 50798 11840 50804 11852
rect 50856 11840 50862 11892
rect 51994 11840 52000 11892
rect 52052 11880 52058 11892
rect 52052 11852 52408 11880
rect 52052 11840 52058 11852
rect 48869 11815 48927 11821
rect 48869 11812 48881 11815
rect 47872 11784 48881 11812
rect 48869 11781 48881 11784
rect 48915 11781 48927 11815
rect 48869 11775 48927 11781
rect 48958 11772 48964 11824
rect 49016 11812 49022 11824
rect 49016 11784 51028 11812
rect 49016 11772 49022 11784
rect 45741 11747 45799 11753
rect 45741 11713 45753 11747
rect 45787 11713 45799 11747
rect 45741 11707 45799 11713
rect 45833 11747 45891 11753
rect 45833 11713 45845 11747
rect 45879 11744 45891 11747
rect 46106 11744 46112 11756
rect 45879 11716 46112 11744
rect 45879 11713 45891 11716
rect 45833 11707 45891 11713
rect 46106 11704 46112 11716
rect 46164 11704 46170 11756
rect 46198 11704 46204 11756
rect 46256 11744 46262 11756
rect 46385 11747 46443 11753
rect 46385 11744 46397 11747
rect 46256 11716 46397 11744
rect 46256 11704 46262 11716
rect 46385 11713 46397 11716
rect 46431 11713 46443 11747
rect 46385 11707 46443 11713
rect 46845 11747 46903 11753
rect 46845 11713 46857 11747
rect 46891 11744 46903 11747
rect 48590 11744 48596 11756
rect 46891 11716 48360 11744
rect 48551 11716 48596 11744
rect 46891 11713 46903 11716
rect 46845 11707 46903 11713
rect 33796 11648 34836 11676
rect 34885 11679 34943 11685
rect 34885 11645 34897 11679
rect 34931 11676 34943 11679
rect 35345 11679 35403 11685
rect 35345 11676 35357 11679
rect 34931 11648 35357 11676
rect 34931 11645 34943 11648
rect 34885 11639 34943 11645
rect 35345 11645 35357 11648
rect 35391 11645 35403 11679
rect 35897 11679 35955 11685
rect 35897 11676 35909 11679
rect 35345 11639 35403 11645
rect 35452 11648 35909 11676
rect 32490 11608 32496 11620
rect 32324 11580 32496 11608
rect 31352 11568 31358 11580
rect 32490 11568 32496 11580
rect 32548 11568 32554 11620
rect 35452 11608 35480 11648
rect 35897 11645 35909 11648
rect 35943 11645 35955 11679
rect 36096 11676 36124 11704
rect 36998 11676 37004 11688
rect 36096 11648 37004 11676
rect 35897 11639 35955 11645
rect 36998 11636 37004 11648
rect 37056 11676 37062 11688
rect 37056 11648 37504 11676
rect 37056 11636 37062 11648
rect 32600 11580 35480 11608
rect 35713 11611 35771 11617
rect 27341 11543 27399 11549
rect 27341 11540 27353 11543
rect 27304 11512 27353 11540
rect 27304 11500 27310 11512
rect 27341 11509 27353 11512
rect 27387 11509 27399 11543
rect 27341 11503 27399 11509
rect 27522 11500 27528 11552
rect 27580 11540 27586 11552
rect 28077 11543 28135 11549
rect 28077 11540 28089 11543
rect 27580 11512 28089 11540
rect 27580 11500 27586 11512
rect 28077 11509 28089 11512
rect 28123 11509 28135 11543
rect 29822 11540 29828 11552
rect 29783 11512 29828 11540
rect 28077 11503 28135 11509
rect 29822 11500 29828 11512
rect 29880 11500 29886 11552
rect 31662 11500 31668 11552
rect 31720 11540 31726 11552
rect 32600 11540 32628 11580
rect 35713 11577 35725 11611
rect 35759 11608 35771 11611
rect 35759 11580 36768 11608
rect 35759 11577 35771 11580
rect 35713 11571 35771 11577
rect 36740 11552 36768 11580
rect 31720 11512 32628 11540
rect 31720 11500 31726 11512
rect 33226 11500 33232 11552
rect 33284 11540 33290 11552
rect 33962 11540 33968 11552
rect 33284 11512 33968 11540
rect 33284 11500 33290 11512
rect 33962 11500 33968 11512
rect 34020 11500 34026 11552
rect 34793 11543 34851 11549
rect 34793 11509 34805 11543
rect 34839 11540 34851 11543
rect 35342 11540 35348 11552
rect 34839 11512 35348 11540
rect 34839 11509 34851 11512
rect 34793 11503 34851 11509
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 35805 11543 35863 11549
rect 35805 11509 35817 11543
rect 35851 11540 35863 11543
rect 36078 11540 36084 11552
rect 35851 11512 36084 11540
rect 35851 11509 35863 11512
rect 35805 11503 35863 11509
rect 36078 11500 36084 11512
rect 36136 11500 36142 11552
rect 36722 11540 36728 11552
rect 36683 11512 36728 11540
rect 36722 11500 36728 11512
rect 36780 11500 36786 11552
rect 37476 11540 37504 11648
rect 37734 11636 37740 11688
rect 37792 11676 37798 11688
rect 37829 11679 37887 11685
rect 37829 11676 37841 11679
rect 37792 11648 37841 11676
rect 37792 11636 37798 11648
rect 37829 11645 37841 11648
rect 37875 11645 37887 11679
rect 37829 11639 37887 11645
rect 38013 11679 38071 11685
rect 38013 11645 38025 11679
rect 38059 11676 38071 11679
rect 38470 11676 38476 11688
rect 38059 11648 38476 11676
rect 38059 11645 38071 11648
rect 38013 11639 38071 11645
rect 38470 11636 38476 11648
rect 38528 11636 38534 11688
rect 41785 11679 41843 11685
rect 41785 11645 41797 11679
rect 41831 11676 41843 11679
rect 42794 11676 42800 11688
rect 41831 11648 42800 11676
rect 41831 11645 41843 11648
rect 41785 11639 41843 11645
rect 42794 11636 42800 11648
rect 42852 11636 42858 11688
rect 43990 11636 43996 11688
rect 44048 11676 44054 11688
rect 44821 11679 44879 11685
rect 44821 11676 44833 11679
rect 44048 11648 44833 11676
rect 44048 11636 44054 11648
rect 44821 11645 44833 11648
rect 44867 11676 44879 11679
rect 46661 11679 46719 11685
rect 46661 11676 46673 11679
rect 44867 11648 46673 11676
rect 44867 11645 44879 11648
rect 44821 11639 44879 11645
rect 46661 11645 46673 11648
rect 46707 11645 46719 11679
rect 46661 11639 46719 11645
rect 37550 11568 37556 11620
rect 37608 11608 37614 11620
rect 38930 11608 38936 11620
rect 37608 11580 38936 11608
rect 37608 11568 37614 11580
rect 38930 11568 38936 11580
rect 38988 11568 38994 11620
rect 43257 11611 43315 11617
rect 43257 11577 43269 11611
rect 43303 11608 43315 11611
rect 45094 11608 45100 11620
rect 43303 11580 45100 11608
rect 43303 11577 43315 11580
rect 43257 11571 43315 11577
rect 45094 11568 45100 11580
rect 45152 11608 45158 11620
rect 45646 11608 45652 11620
rect 45152 11580 45508 11608
rect 45607 11580 45652 11608
rect 45152 11568 45158 11580
rect 37918 11540 37924 11552
rect 37476 11512 37924 11540
rect 37918 11500 37924 11512
rect 37976 11500 37982 11552
rect 39206 11540 39212 11552
rect 39167 11512 39212 11540
rect 39206 11500 39212 11512
rect 39264 11500 39270 11552
rect 40221 11543 40279 11549
rect 40221 11509 40233 11543
rect 40267 11540 40279 11543
rect 40402 11540 40408 11552
rect 40267 11512 40408 11540
rect 40267 11509 40279 11512
rect 40221 11503 40279 11509
rect 40402 11500 40408 11512
rect 40460 11500 40466 11552
rect 43346 11500 43352 11552
rect 43404 11540 43410 11552
rect 45480 11540 45508 11580
rect 45646 11568 45652 11580
rect 45704 11568 45710 11620
rect 47765 11611 47823 11617
rect 47765 11608 47777 11611
rect 45940 11580 47777 11608
rect 45940 11540 45968 11580
rect 47765 11577 47777 11580
rect 47811 11577 47823 11611
rect 47765 11571 47823 11577
rect 43404 11512 43449 11540
rect 45480 11512 45968 11540
rect 46523 11543 46581 11549
rect 43404 11500 43410 11512
rect 46523 11509 46535 11543
rect 46569 11540 46581 11543
rect 46750 11540 46756 11552
rect 46569 11512 46756 11540
rect 46569 11509 46581 11512
rect 46523 11503 46581 11509
rect 46750 11500 46756 11512
rect 46808 11500 46814 11552
rect 48332 11540 48360 11716
rect 48590 11704 48596 11716
rect 48648 11704 48654 11756
rect 48682 11704 48688 11756
rect 48740 11744 48746 11756
rect 49421 11747 49479 11753
rect 49421 11744 49433 11747
rect 48740 11716 49433 11744
rect 48740 11704 48746 11716
rect 49421 11713 49433 11716
rect 49467 11713 49479 11747
rect 49421 11707 49479 11713
rect 50798 11747 50856 11753
rect 50798 11713 50810 11747
rect 50844 11744 50856 11747
rect 50844 11716 50948 11744
rect 50844 11713 50856 11716
rect 50798 11707 50856 11713
rect 48501 11679 48559 11685
rect 48501 11645 48513 11679
rect 48547 11645 48559 11679
rect 48501 11639 48559 11645
rect 48516 11608 48544 11639
rect 48774 11636 48780 11688
rect 48832 11676 48838 11688
rect 48961 11679 49019 11685
rect 48961 11676 48973 11679
rect 48832 11648 48973 11676
rect 48832 11636 48838 11648
rect 48961 11645 48973 11648
rect 49007 11676 49019 11679
rect 49142 11676 49148 11688
rect 49007 11648 49148 11676
rect 49007 11645 49019 11648
rect 48961 11639 49019 11645
rect 49142 11636 49148 11648
rect 49200 11636 49206 11688
rect 49510 11676 49516 11688
rect 49471 11648 49516 11676
rect 49510 11636 49516 11648
rect 49568 11636 49574 11688
rect 50920 11608 50948 11716
rect 51000 11676 51028 11784
rect 51074 11772 51080 11824
rect 51132 11812 51138 11824
rect 51132 11784 52316 11812
rect 51132 11772 51138 11784
rect 51261 11747 51319 11753
rect 51261 11713 51273 11747
rect 51307 11744 51319 11747
rect 51997 11747 52055 11753
rect 51997 11745 52009 11747
rect 51920 11744 52009 11745
rect 51307 11716 51764 11744
rect 51307 11713 51319 11716
rect 51261 11707 51319 11713
rect 51169 11679 51227 11685
rect 51169 11676 51181 11679
rect 51000 11648 51181 11676
rect 51169 11645 51181 11648
rect 51215 11676 51227 11679
rect 51626 11676 51632 11688
rect 51215 11648 51632 11676
rect 51215 11645 51227 11648
rect 51169 11639 51227 11645
rect 51626 11636 51632 11648
rect 51684 11636 51690 11688
rect 51736 11685 51764 11716
rect 51828 11717 52009 11744
rect 51828 11716 51948 11717
rect 51721 11679 51779 11685
rect 51721 11645 51733 11679
rect 51767 11645 51779 11679
rect 51721 11639 51779 11645
rect 51350 11608 51356 11620
rect 48516 11580 48820 11608
rect 50920 11580 51356 11608
rect 48792 11552 48820 11580
rect 51350 11568 51356 11580
rect 51408 11568 51414 11620
rect 48498 11540 48504 11552
rect 48332 11512 48504 11540
rect 48498 11500 48504 11512
rect 48556 11500 48562 11552
rect 48774 11500 48780 11552
rect 48832 11500 48838 11552
rect 49418 11540 49424 11552
rect 49379 11512 49424 11540
rect 49418 11500 49424 11512
rect 49476 11500 49482 11552
rect 51368 11540 51396 11568
rect 51718 11540 51724 11552
rect 51368 11512 51724 11540
rect 51718 11500 51724 11512
rect 51776 11500 51782 11552
rect 51828 11540 51856 11716
rect 51997 11713 52009 11717
rect 52043 11713 52055 11747
rect 51997 11707 52055 11713
rect 52089 11747 52147 11753
rect 52089 11713 52101 11747
rect 52135 11713 52147 11747
rect 52089 11707 52147 11713
rect 52181 11747 52239 11753
rect 52181 11713 52193 11747
rect 52227 11745 52239 11747
rect 52288 11745 52316 11784
rect 52380 11756 52408 11852
rect 52546 11840 52552 11892
rect 52604 11880 52610 11892
rect 53929 11883 53987 11889
rect 53929 11880 53941 11883
rect 52604 11852 53941 11880
rect 52604 11840 52610 11852
rect 53929 11849 53941 11852
rect 53975 11880 53987 11883
rect 54202 11880 54208 11892
rect 53975 11852 54208 11880
rect 53975 11849 53987 11852
rect 53929 11843 53987 11849
rect 54202 11840 54208 11852
rect 54260 11840 54266 11892
rect 54297 11883 54355 11889
rect 54297 11849 54309 11883
rect 54343 11880 54355 11883
rect 55674 11880 55680 11892
rect 54343 11852 55680 11880
rect 54343 11849 54355 11852
rect 54297 11843 54355 11849
rect 55674 11840 55680 11852
rect 55732 11840 55738 11892
rect 55950 11880 55956 11892
rect 55911 11852 55956 11880
rect 55950 11840 55956 11852
rect 56008 11840 56014 11892
rect 53190 11772 53196 11824
rect 53248 11812 53254 11824
rect 54478 11812 54484 11824
rect 53248 11784 54484 11812
rect 53248 11772 53254 11784
rect 54478 11772 54484 11784
rect 54536 11812 54542 11824
rect 54536 11784 55260 11812
rect 54536 11772 54542 11784
rect 52227 11717 52316 11745
rect 52227 11713 52239 11717
rect 52181 11707 52239 11713
rect 52104 11620 52132 11707
rect 52362 11704 52368 11756
rect 52420 11744 52426 11756
rect 52420 11716 52513 11744
rect 52420 11704 52426 11716
rect 53558 11704 53564 11756
rect 53616 11744 53622 11756
rect 53837 11747 53895 11753
rect 53837 11744 53849 11747
rect 53616 11716 53849 11744
rect 53616 11704 53622 11716
rect 53837 11713 53849 11716
rect 53883 11713 53895 11747
rect 54110 11744 54116 11756
rect 54023 11716 54116 11744
rect 53837 11707 53895 11713
rect 54110 11704 54116 11716
rect 54168 11704 54174 11756
rect 54570 11704 54576 11756
rect 54628 11744 54634 11756
rect 54849 11747 54907 11753
rect 54849 11744 54861 11747
rect 54628 11716 54861 11744
rect 54628 11704 54634 11716
rect 54849 11713 54861 11716
rect 54895 11713 54907 11747
rect 55030 11744 55036 11756
rect 54991 11716 55036 11744
rect 54849 11707 54907 11713
rect 55030 11704 55036 11716
rect 55088 11704 55094 11756
rect 55232 11744 55260 11784
rect 55490 11772 55496 11824
rect 55548 11812 55554 11824
rect 55585 11815 55643 11821
rect 55585 11812 55597 11815
rect 55548 11784 55597 11812
rect 55548 11772 55554 11784
rect 55585 11781 55597 11784
rect 55631 11781 55643 11815
rect 55585 11775 55643 11781
rect 55766 11772 55772 11824
rect 55824 11821 55830 11824
rect 55824 11815 55843 11821
rect 55831 11781 55843 11815
rect 55824 11775 55843 11781
rect 55824 11772 55830 11775
rect 56965 11747 57023 11753
rect 56965 11744 56977 11747
rect 55232 11716 56977 11744
rect 56965 11713 56977 11716
rect 57011 11713 57023 11747
rect 56965 11707 57023 11713
rect 53374 11636 53380 11688
rect 53432 11676 53438 11688
rect 54128 11676 54156 11704
rect 53432 11648 54156 11676
rect 53432 11636 53438 11648
rect 54202 11636 54208 11688
rect 54260 11676 54266 11688
rect 55048 11676 55076 11704
rect 54260 11648 55076 11676
rect 54260 11636 54266 11648
rect 52086 11568 52092 11620
rect 52144 11568 52150 11620
rect 53282 11608 53288 11620
rect 52196 11580 53288 11608
rect 52196 11540 52224 11580
rect 53282 11568 53288 11580
rect 53340 11568 53346 11620
rect 54846 11608 54852 11620
rect 54807 11580 54852 11608
rect 54846 11568 54852 11580
rect 54904 11568 54910 11620
rect 55048 11608 55076 11648
rect 55048 11580 55812 11608
rect 51828 11512 52224 11540
rect 52730 11500 52736 11552
rect 52788 11540 52794 11552
rect 52917 11543 52975 11549
rect 52917 11540 52929 11543
rect 52788 11512 52929 11540
rect 52788 11500 52794 11512
rect 52917 11509 52929 11512
rect 52963 11540 52975 11543
rect 55674 11540 55680 11552
rect 52963 11512 55680 11540
rect 52963 11509 52975 11512
rect 52917 11503 52975 11509
rect 55674 11500 55680 11512
rect 55732 11500 55738 11552
rect 55784 11549 55812 11580
rect 55769 11543 55827 11549
rect 55769 11509 55781 11543
rect 55815 11509 55827 11543
rect 55769 11503 55827 11509
rect 56505 11543 56563 11549
rect 56505 11509 56517 11543
rect 56551 11540 56563 11543
rect 57422 11540 57428 11552
rect 56551 11512 57428 11540
rect 56551 11509 56563 11512
rect 56505 11503 56563 11509
rect 57422 11500 57428 11512
rect 57480 11540 57486 11552
rect 57882 11540 57888 11552
rect 57480 11512 57888 11540
rect 57480 11500 57486 11512
rect 57882 11500 57888 11512
rect 57940 11500 57946 11552
rect 58161 11543 58219 11549
rect 58161 11509 58173 11543
rect 58207 11540 58219 11543
rect 58250 11540 58256 11552
rect 58207 11512 58256 11540
rect 58207 11509 58219 11512
rect 58161 11503 58219 11509
rect 58250 11500 58256 11512
rect 58308 11500 58314 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 25593 11339 25651 11345
rect 25593 11305 25605 11339
rect 25639 11336 25651 11339
rect 26050 11336 26056 11348
rect 25639 11308 26056 11336
rect 25639 11305 25651 11308
rect 25593 11299 25651 11305
rect 26050 11296 26056 11308
rect 26108 11296 26114 11348
rect 27430 11336 27436 11348
rect 27391 11308 27436 11336
rect 27430 11296 27436 11308
rect 27488 11296 27494 11348
rect 28258 11336 28264 11348
rect 28219 11308 28264 11336
rect 28258 11296 28264 11308
rect 28316 11336 28322 11348
rect 28810 11336 28816 11348
rect 28316 11308 28816 11336
rect 28316 11296 28322 11308
rect 28810 11296 28816 11308
rect 28868 11296 28874 11348
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 29825 11339 29883 11345
rect 29825 11336 29837 11339
rect 29052 11308 29837 11336
rect 29052 11296 29058 11308
rect 29825 11305 29837 11308
rect 29871 11305 29883 11339
rect 29825 11299 29883 11305
rect 30561 11339 30619 11345
rect 30561 11305 30573 11339
rect 30607 11336 30619 11339
rect 30650 11336 30656 11348
rect 30607 11308 30656 11336
rect 30607 11305 30619 11308
rect 30561 11299 30619 11305
rect 25682 11228 25688 11280
rect 25740 11268 25746 11280
rect 26329 11271 26387 11277
rect 26329 11268 26341 11271
rect 25740 11240 26341 11268
rect 25740 11228 25746 11240
rect 26329 11237 26341 11240
rect 26375 11237 26387 11271
rect 26329 11231 26387 11237
rect 27338 11228 27344 11280
rect 27396 11268 27402 11280
rect 28902 11268 28908 11280
rect 27396 11240 28908 11268
rect 27396 11228 27402 11240
rect 28902 11228 28908 11240
rect 28960 11268 28966 11280
rect 29454 11268 29460 11280
rect 28960 11240 29460 11268
rect 28960 11228 28966 11240
rect 29454 11228 29460 11240
rect 29512 11228 29518 11280
rect 29840 11268 29868 11299
rect 30650 11296 30656 11308
rect 30708 11296 30714 11348
rect 32125 11339 32183 11345
rect 32125 11305 32137 11339
rect 32171 11336 32183 11339
rect 32306 11336 32312 11348
rect 32171 11308 32312 11336
rect 32171 11305 32183 11308
rect 32125 11299 32183 11305
rect 32306 11296 32312 11308
rect 32364 11296 32370 11348
rect 32950 11336 32956 11348
rect 32911 11308 32956 11336
rect 32950 11296 32956 11308
rect 33008 11296 33014 11348
rect 33778 11296 33784 11348
rect 33836 11336 33842 11348
rect 33873 11339 33931 11345
rect 33873 11336 33885 11339
rect 33836 11308 33885 11336
rect 33836 11296 33842 11308
rect 33873 11305 33885 11308
rect 33919 11336 33931 11339
rect 33962 11336 33968 11348
rect 33919 11308 33968 11336
rect 33919 11305 33931 11308
rect 33873 11299 33931 11305
rect 33962 11296 33968 11308
rect 34020 11296 34026 11348
rect 34333 11339 34391 11345
rect 34333 11305 34345 11339
rect 34379 11336 34391 11339
rect 35618 11336 35624 11348
rect 34379 11308 35624 11336
rect 34379 11305 34391 11308
rect 34333 11299 34391 11305
rect 35618 11296 35624 11308
rect 35676 11296 35682 11348
rect 35894 11296 35900 11348
rect 35952 11336 35958 11348
rect 36081 11339 36139 11345
rect 36081 11336 36093 11339
rect 35952 11308 36093 11336
rect 35952 11296 35958 11308
rect 36081 11305 36093 11308
rect 36127 11336 36139 11339
rect 36354 11336 36360 11348
rect 36127 11308 36360 11336
rect 36127 11305 36139 11308
rect 36081 11299 36139 11305
rect 36354 11296 36360 11308
rect 36412 11296 36418 11348
rect 37734 11336 37740 11348
rect 37695 11308 37740 11336
rect 37734 11296 37740 11308
rect 37792 11296 37798 11348
rect 37918 11296 37924 11348
rect 37976 11336 37982 11348
rect 38562 11336 38568 11348
rect 37976 11308 38568 11336
rect 37976 11296 37982 11308
rect 38562 11296 38568 11308
rect 38620 11336 38626 11348
rect 38657 11339 38715 11345
rect 38657 11336 38669 11339
rect 38620 11308 38669 11336
rect 38620 11296 38626 11308
rect 38657 11305 38669 11308
rect 38703 11305 38715 11339
rect 40770 11336 40776 11348
rect 40731 11308 40776 11336
rect 38657 11299 38715 11305
rect 40770 11296 40776 11308
rect 40828 11296 40834 11348
rect 42334 11336 42340 11348
rect 42295 11308 42340 11336
rect 42334 11296 42340 11308
rect 42392 11296 42398 11348
rect 43073 11339 43131 11345
rect 43073 11305 43085 11339
rect 43119 11336 43131 11339
rect 43346 11336 43352 11348
rect 43119 11308 43352 11336
rect 43119 11305 43131 11308
rect 43073 11299 43131 11305
rect 43346 11296 43352 11308
rect 43404 11296 43410 11348
rect 43990 11336 43996 11348
rect 43951 11308 43996 11336
rect 43990 11296 43996 11308
rect 44048 11296 44054 11348
rect 46385 11339 46443 11345
rect 46385 11336 46397 11339
rect 44146 11308 46397 11336
rect 33502 11268 33508 11280
rect 29840 11240 33508 11268
rect 33502 11228 33508 11240
rect 33560 11268 33566 11280
rect 33560 11240 33824 11268
rect 33560 11228 33566 11240
rect 24581 11203 24639 11209
rect 24581 11169 24593 11203
rect 24627 11200 24639 11203
rect 27356 11200 27384 11228
rect 24627 11172 27384 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 27890 11160 27896 11212
rect 27948 11200 27954 11212
rect 30282 11200 30288 11212
rect 27948 11172 30288 11200
rect 27948 11160 27954 11172
rect 30282 11160 30288 11172
rect 30340 11160 30346 11212
rect 30837 11203 30895 11209
rect 30837 11169 30849 11203
rect 30883 11200 30895 11203
rect 31662 11200 31668 11212
rect 30883 11172 31668 11200
rect 30883 11169 30895 11172
rect 30837 11163 30895 11169
rect 31662 11160 31668 11172
rect 31720 11160 31726 11212
rect 33042 11200 33048 11212
rect 32232 11172 33048 11200
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 23842 11024 23848 11076
rect 23900 11064 23906 11076
rect 24780 11064 24808 11095
rect 25038 11092 25044 11144
rect 25096 11132 25102 11144
rect 25409 11135 25467 11141
rect 25409 11132 25421 11135
rect 25096 11104 25421 11132
rect 25096 11092 25102 11104
rect 25409 11101 25421 11104
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 25593 11135 25651 11141
rect 25593 11101 25605 11135
rect 25639 11132 25651 11135
rect 25958 11132 25964 11144
rect 25639 11104 25964 11132
rect 25639 11101 25651 11104
rect 25593 11095 25651 11101
rect 23900 11036 24808 11064
rect 25424 11064 25452 11095
rect 25958 11092 25964 11104
rect 26016 11092 26022 11144
rect 27801 11135 27859 11141
rect 27801 11101 27813 11135
rect 27847 11132 27859 11135
rect 28166 11132 28172 11144
rect 27847 11104 28172 11132
rect 27847 11101 27859 11104
rect 27801 11095 27859 11101
rect 28166 11092 28172 11104
rect 28224 11092 28230 11144
rect 28350 11092 28356 11144
rect 28408 11132 28414 11144
rect 28445 11135 28503 11141
rect 28445 11132 28457 11135
rect 28408 11104 28457 11132
rect 28408 11092 28414 11104
rect 28445 11101 28457 11104
rect 28491 11101 28503 11135
rect 28629 11135 28687 11141
rect 28629 11132 28641 11135
rect 28445 11095 28503 11101
rect 28552 11104 28641 11132
rect 26142 11064 26148 11076
rect 25424 11036 26148 11064
rect 23900 11024 23906 11036
rect 26142 11024 26148 11036
rect 26200 11024 26206 11076
rect 27614 11064 27620 11076
rect 27575 11036 27620 11064
rect 27614 11024 27620 11036
rect 27672 11024 27678 11076
rect 28258 11024 28264 11076
rect 28316 11064 28322 11076
rect 28552 11064 28580 11104
rect 28629 11101 28641 11104
rect 28675 11101 28687 11135
rect 28629 11095 28687 11101
rect 28721 11135 28779 11141
rect 28721 11101 28733 11135
rect 28767 11134 28779 11135
rect 28767 11106 28856 11134
rect 28767 11101 28779 11106
rect 28721 11095 28779 11101
rect 28316 11036 28580 11064
rect 28828 11064 28856 11106
rect 28902 11092 28908 11144
rect 28960 11132 28966 11144
rect 29733 11135 29791 11141
rect 28960 11126 29684 11132
rect 29733 11126 29745 11135
rect 28960 11104 29745 11126
rect 28960 11092 28966 11104
rect 29454 11064 29460 11076
rect 28828 11036 29460 11064
rect 28316 11024 28322 11036
rect 29454 11024 29460 11036
rect 29512 11024 29518 11076
rect 29564 11064 29592 11104
rect 29656 11101 29745 11104
rect 29779 11101 29791 11135
rect 29656 11098 29791 11101
rect 29733 11095 29791 11098
rect 29914 11092 29920 11144
rect 29972 11132 29978 11144
rect 29972 11104 30017 11132
rect 29972 11092 29978 11104
rect 30558 11092 30564 11144
rect 30616 11132 30622 11144
rect 30745 11135 30803 11141
rect 30745 11132 30757 11135
rect 30616 11104 30757 11132
rect 30616 11092 30622 11104
rect 30745 11101 30757 11104
rect 30791 11101 30803 11135
rect 30745 11095 30803 11101
rect 30926 11092 30932 11144
rect 30984 11132 30990 11144
rect 31057 11135 31115 11141
rect 30984 11104 31029 11132
rect 30984 11092 30990 11104
rect 31057 11101 31069 11135
rect 31103 11132 31115 11135
rect 31202 11132 31208 11144
rect 31103 11104 31208 11132
rect 31103 11101 31115 11104
rect 31057 11095 31115 11101
rect 31202 11092 31208 11104
rect 31260 11092 31266 11144
rect 32030 11132 32036 11144
rect 31991 11104 32036 11132
rect 32030 11092 32036 11104
rect 32088 11092 32094 11144
rect 32232 11141 32260 11172
rect 33042 11160 33048 11172
rect 33100 11160 33106 11212
rect 33796 11141 33824 11240
rect 34882 11228 34888 11280
rect 34940 11268 34946 11280
rect 35802 11268 35808 11280
rect 34940 11240 35808 11268
rect 34940 11228 34946 11240
rect 35802 11228 35808 11240
rect 35860 11228 35866 11280
rect 36538 11268 36544 11280
rect 36499 11240 36544 11268
rect 36538 11228 36544 11240
rect 36596 11228 36602 11280
rect 37274 11228 37280 11280
rect 37332 11268 37338 11280
rect 38102 11268 38108 11280
rect 37332 11240 38108 11268
rect 37332 11228 37338 11240
rect 38102 11228 38108 11240
rect 38160 11228 38166 11280
rect 39390 11228 39396 11280
rect 39448 11268 39454 11280
rect 41233 11271 41291 11277
rect 41233 11268 41245 11271
rect 39448 11240 41245 11268
rect 39448 11228 39454 11240
rect 41233 11237 41245 11240
rect 41279 11237 41291 11271
rect 41233 11231 41291 11237
rect 43714 11228 43720 11280
rect 43772 11268 43778 11280
rect 44146 11268 44174 11308
rect 46385 11305 46397 11308
rect 46431 11305 46443 11339
rect 46385 11299 46443 11305
rect 46934 11296 46940 11348
rect 46992 11336 46998 11348
rect 47762 11336 47768 11348
rect 46992 11308 47768 11336
rect 46992 11296 46998 11308
rect 47762 11296 47768 11308
rect 47820 11296 47826 11348
rect 48317 11339 48375 11345
rect 48317 11305 48329 11339
rect 48363 11336 48375 11339
rect 48682 11336 48688 11348
rect 48363 11308 48688 11336
rect 48363 11305 48375 11308
rect 48317 11299 48375 11305
rect 48682 11296 48688 11308
rect 48740 11296 48746 11348
rect 49050 11296 49056 11348
rect 49108 11336 49114 11348
rect 49605 11339 49663 11345
rect 49605 11336 49617 11339
rect 49108 11308 49617 11336
rect 49108 11296 49114 11308
rect 49605 11305 49617 11308
rect 49651 11336 49663 11339
rect 49651 11308 50844 11336
rect 49651 11305 49663 11308
rect 49605 11299 49663 11305
rect 43772 11240 44174 11268
rect 43772 11228 43778 11240
rect 45094 11228 45100 11280
rect 45152 11228 45158 11280
rect 45922 11228 45928 11280
rect 45980 11268 45986 11280
rect 47210 11268 47216 11280
rect 45980 11240 47216 11268
rect 45980 11228 45986 11240
rect 47210 11228 47216 11240
rect 47268 11228 47274 11280
rect 50706 11228 50712 11280
rect 50764 11228 50770 11280
rect 35618 11160 35624 11212
rect 35676 11200 35682 11212
rect 35676 11172 37688 11200
rect 35676 11160 35682 11172
rect 32217 11135 32275 11141
rect 32217 11101 32229 11135
rect 32263 11101 32275 11135
rect 33781 11135 33839 11141
rect 32217 11095 32275 11101
rect 32324 11119 32720 11132
rect 32324 11113 32735 11119
rect 32324 11104 32689 11113
rect 29822 11064 29828 11076
rect 29564 11036 29828 11064
rect 29822 11024 29828 11036
rect 29880 11064 29886 11076
rect 29880 11036 31340 11064
rect 29880 11024 29886 11036
rect 25682 10956 25688 11008
rect 25740 10996 25746 11008
rect 26878 10996 26884 11008
rect 25740 10968 26884 10996
rect 25740 10956 25746 10968
rect 26878 10956 26884 10968
rect 26936 10956 26942 11008
rect 27246 10956 27252 11008
rect 27304 10996 27310 11008
rect 31202 10996 31208 11008
rect 27304 10968 31208 10996
rect 27304 10956 27310 10968
rect 31202 10956 31208 10968
rect 31260 10956 31266 11008
rect 31312 10996 31340 11036
rect 31386 11024 31392 11076
rect 31444 11064 31450 11076
rect 32324 11064 32352 11104
rect 32677 11079 32689 11104
rect 32723 11079 32735 11113
rect 33781 11101 33793 11135
rect 33827 11101 33839 11135
rect 33781 11095 33839 11101
rect 34149 11135 34207 11141
rect 34149 11101 34161 11135
rect 34195 11132 34207 11135
rect 34422 11132 34428 11144
rect 34195 11104 34428 11132
rect 34195 11101 34207 11104
rect 34149 11095 34207 11101
rect 34422 11092 34428 11104
rect 34480 11092 34486 11144
rect 35526 11092 35532 11144
rect 35584 11132 35590 11144
rect 36814 11132 36820 11144
rect 35584 11104 35629 11132
rect 36775 11104 36820 11132
rect 35584 11092 35590 11104
rect 36814 11092 36820 11104
rect 36872 11092 36878 11144
rect 37182 11092 37188 11144
rect 37240 11132 37246 11144
rect 37277 11135 37335 11141
rect 37277 11132 37289 11135
rect 37240 11104 37289 11132
rect 37240 11092 37246 11104
rect 37277 11101 37289 11104
rect 37323 11101 37335 11135
rect 37550 11132 37556 11144
rect 37511 11104 37556 11132
rect 37277 11095 37335 11101
rect 37550 11092 37556 11104
rect 37608 11092 37614 11144
rect 37660 11132 37688 11172
rect 38654 11160 38660 11212
rect 38712 11200 38718 11212
rect 40129 11203 40187 11209
rect 40129 11200 40141 11203
rect 38712 11172 40141 11200
rect 38712 11160 38718 11172
rect 40129 11169 40141 11172
rect 40175 11169 40187 11203
rect 40129 11163 40187 11169
rect 42702 11160 42708 11212
rect 42760 11200 42766 11212
rect 43162 11200 43168 11212
rect 42760 11172 43168 11200
rect 42760 11160 42766 11172
rect 43162 11160 43168 11172
rect 43220 11200 43226 11212
rect 43220 11172 43576 11200
rect 43220 11160 43226 11172
rect 38841 11135 38899 11141
rect 38841 11132 38853 11135
rect 37660 11104 38853 11132
rect 38841 11101 38853 11104
rect 38887 11132 38899 11135
rect 39022 11132 39028 11144
rect 38887 11104 39028 11132
rect 38887 11101 38899 11104
rect 38841 11095 38899 11101
rect 39022 11092 39028 11104
rect 39080 11092 39086 11144
rect 40402 11132 40408 11144
rect 40363 11104 40408 11132
rect 40402 11092 40408 11104
rect 40460 11092 40466 11144
rect 42610 11092 42616 11144
rect 42668 11132 42674 11144
rect 43548 11141 43576 11172
rect 42889 11135 42947 11141
rect 42889 11132 42901 11135
rect 42668 11104 42901 11132
rect 42668 11092 42674 11104
rect 42889 11101 42901 11104
rect 42935 11101 42947 11135
rect 42889 11095 42947 11101
rect 43073 11135 43131 11141
rect 43073 11101 43085 11135
rect 43119 11101 43131 11135
rect 43073 11095 43131 11101
rect 43533 11135 43591 11141
rect 43533 11101 43545 11135
rect 43579 11101 43591 11135
rect 43533 11095 43591 11101
rect 43809 11135 43867 11141
rect 43809 11101 43821 11135
rect 43855 11132 43867 11135
rect 44818 11132 44824 11144
rect 43855 11104 44824 11132
rect 43855 11101 43867 11104
rect 43809 11095 43867 11101
rect 32677 11073 32735 11079
rect 31444 11036 32352 11064
rect 31444 11024 31450 11036
rect 32766 11024 32772 11076
rect 32824 11064 32830 11076
rect 32824 11036 32869 11064
rect 32824 11024 32830 11036
rect 32950 11024 32956 11076
rect 33008 11064 33014 11076
rect 33008 11036 33053 11064
rect 33008 11024 33014 11036
rect 34238 11024 34244 11076
rect 34296 11064 34302 11076
rect 36541 11067 36599 11073
rect 36541 11064 36553 11067
rect 34296 11036 36553 11064
rect 34296 11024 34302 11036
rect 36541 11033 36553 11036
rect 36587 11033 36599 11067
rect 36541 11027 36599 11033
rect 36725 11067 36783 11073
rect 36725 11033 36737 11067
rect 36771 11064 36783 11067
rect 36906 11064 36912 11076
rect 36771 11036 36912 11064
rect 36771 11033 36783 11036
rect 36725 11027 36783 11033
rect 36906 11024 36912 11036
rect 36964 11024 36970 11076
rect 39301 11067 39359 11073
rect 39301 11064 39313 11067
rect 38626 11036 39313 11064
rect 31662 10996 31668 11008
rect 31312 10968 31668 10996
rect 31662 10956 31668 10968
rect 31720 10956 31726 11008
rect 32968 10996 32996 11024
rect 34885 10999 34943 11005
rect 34885 10996 34897 10999
rect 32968 10968 34897 10996
rect 34885 10965 34897 10968
rect 34931 10996 34943 10999
rect 35434 10996 35440 11008
rect 34931 10968 35440 10996
rect 34931 10965 34943 10968
rect 34885 10959 34943 10965
rect 35434 10956 35440 10968
rect 35492 10956 35498 11008
rect 37366 10996 37372 11008
rect 37327 10968 37372 10996
rect 37366 10956 37372 10968
rect 37424 10996 37430 11008
rect 38626 10996 38654 11036
rect 39301 11033 39313 11036
rect 39347 11033 39359 11067
rect 39301 11027 39359 11033
rect 40218 11024 40224 11076
rect 40276 11064 40282 11076
rect 40313 11067 40371 11073
rect 40313 11064 40325 11067
rect 40276 11036 40325 11064
rect 40276 11024 40282 11036
rect 40313 11033 40325 11036
rect 40359 11033 40371 11067
rect 40313 11027 40371 11033
rect 41782 10996 41788 11008
rect 37424 10968 38654 10996
rect 41743 10968 41788 10996
rect 37424 10956 37430 10968
rect 41782 10956 41788 10968
rect 41840 10956 41846 11008
rect 43088 10996 43116 11095
rect 44818 11092 44824 11104
rect 44876 11092 44882 11144
rect 45112 11132 45140 11228
rect 45281 11203 45339 11209
rect 45281 11169 45293 11203
rect 45327 11200 45339 11203
rect 45554 11200 45560 11212
rect 45327 11172 45560 11200
rect 45327 11169 45339 11172
rect 45281 11163 45339 11169
rect 45554 11160 45560 11172
rect 45612 11200 45618 11212
rect 47397 11203 47455 11209
rect 47397 11200 47409 11203
rect 45612 11172 47409 11200
rect 45612 11160 45618 11172
rect 47397 11169 47409 11172
rect 47443 11169 47455 11203
rect 47397 11163 47455 11169
rect 47486 11160 47492 11212
rect 47544 11200 47550 11212
rect 48961 11203 49019 11209
rect 48961 11200 48973 11203
rect 47544 11172 47589 11200
rect 47688 11172 48973 11200
rect 47544 11160 47550 11172
rect 45181 11135 45239 11141
rect 45181 11132 45193 11135
rect 45112 11104 45193 11132
rect 45181 11101 45193 11104
rect 45227 11101 45239 11135
rect 47302 11132 47308 11144
rect 47263 11104 47308 11132
rect 45181 11095 45239 11101
rect 47302 11092 47308 11104
rect 47360 11092 47366 11144
rect 47578 11132 47584 11144
rect 47539 11104 47584 11132
rect 47578 11092 47584 11104
rect 47636 11092 47642 11144
rect 43162 11024 43168 11076
rect 43220 11064 43226 11076
rect 43625 11067 43683 11073
rect 43625 11064 43637 11067
rect 43220 11036 43637 11064
rect 43220 11024 43226 11036
rect 43625 11033 43637 11036
rect 43671 11033 43683 11067
rect 44542 11064 44548 11076
rect 44455 11036 44548 11064
rect 43625 11027 43683 11033
rect 44542 11024 44548 11036
rect 44600 11064 44606 11076
rect 45738 11064 45744 11076
rect 44600 11036 45744 11064
rect 44600 11024 44606 11036
rect 45738 11024 45744 11036
rect 45796 11024 45802 11076
rect 47394 11024 47400 11076
rect 47452 11064 47458 11076
rect 47688 11064 47716 11172
rect 48961 11169 48973 11172
rect 49007 11169 49019 11203
rect 50724 11200 50752 11228
rect 48961 11163 49019 11169
rect 50356 11172 50752 11200
rect 47762 11092 47768 11144
rect 47820 11092 47826 11144
rect 48314 11092 48320 11144
rect 48372 11132 48378 11144
rect 48498 11132 48504 11144
rect 48372 11104 48417 11132
rect 48459 11104 48504 11132
rect 48372 11092 48378 11104
rect 48498 11092 48504 11104
rect 48556 11092 48562 11144
rect 48774 11092 48780 11144
rect 48832 11132 48838 11144
rect 49970 11132 49976 11144
rect 48832 11104 49976 11132
rect 48832 11092 48838 11104
rect 49970 11092 49976 11104
rect 50028 11132 50034 11144
rect 50154 11132 50160 11144
rect 50028 11104 50160 11132
rect 50028 11092 50034 11104
rect 50154 11092 50160 11104
rect 50212 11092 50218 11144
rect 50356 11141 50384 11172
rect 50341 11135 50399 11141
rect 50341 11101 50353 11135
rect 50387 11101 50399 11135
rect 50522 11132 50528 11144
rect 50483 11104 50528 11132
rect 50341 11095 50399 11101
rect 50522 11092 50528 11104
rect 50580 11092 50586 11144
rect 50617 11135 50675 11141
rect 50617 11101 50629 11135
rect 50663 11101 50675 11135
rect 50617 11095 50675 11101
rect 50709 11135 50767 11141
rect 50709 11101 50721 11135
rect 50755 11132 50767 11135
rect 50816 11132 50844 11308
rect 50890 11296 50896 11348
rect 50948 11336 50954 11348
rect 50985 11339 51043 11345
rect 50985 11336 50997 11339
rect 50948 11308 50997 11336
rect 50948 11296 50954 11308
rect 50985 11305 50997 11308
rect 51031 11305 51043 11339
rect 50985 11299 51043 11305
rect 52178 11296 52184 11348
rect 52236 11336 52242 11348
rect 53009 11339 53067 11345
rect 53009 11336 53021 11339
rect 52236 11308 53021 11336
rect 52236 11296 52242 11308
rect 53009 11305 53021 11308
rect 53055 11336 53067 11339
rect 54202 11336 54208 11348
rect 53055 11308 54208 11336
rect 53055 11305 53067 11308
rect 53009 11299 53067 11305
rect 54202 11296 54208 11308
rect 54260 11296 54266 11348
rect 54294 11296 54300 11348
rect 54352 11336 54358 11348
rect 54389 11339 54447 11345
rect 54389 11336 54401 11339
rect 54352 11308 54401 11336
rect 54352 11296 54358 11308
rect 54389 11305 54401 11308
rect 54435 11305 54447 11339
rect 54389 11299 54447 11305
rect 55766 11296 55772 11348
rect 55824 11336 55830 11348
rect 55861 11339 55919 11345
rect 55861 11336 55873 11339
rect 55824 11308 55873 11336
rect 55824 11296 55830 11308
rect 55861 11305 55873 11308
rect 55907 11305 55919 11339
rect 58066 11336 58072 11348
rect 58027 11308 58072 11336
rect 55861 11299 55919 11305
rect 51074 11228 51080 11280
rect 51132 11268 51138 11280
rect 51721 11271 51779 11277
rect 51721 11268 51733 11271
rect 51132 11240 51733 11268
rect 51132 11228 51138 11240
rect 51721 11237 51733 11240
rect 51767 11237 51779 11271
rect 52825 11271 52883 11277
rect 52825 11268 52837 11271
rect 51721 11231 51779 11237
rect 52196 11240 52837 11268
rect 52089 11203 52147 11209
rect 52089 11169 52101 11203
rect 52135 11200 52147 11203
rect 52196 11200 52224 11240
rect 52825 11237 52837 11240
rect 52871 11237 52883 11271
rect 52825 11231 52883 11237
rect 52135 11172 52224 11200
rect 52135 11169 52147 11172
rect 52089 11163 52147 11169
rect 53742 11160 53748 11212
rect 53800 11200 53806 11212
rect 53929 11203 53987 11209
rect 53929 11200 53941 11203
rect 53800 11172 53941 11200
rect 53800 11160 53806 11172
rect 53929 11169 53941 11172
rect 53975 11169 53987 11203
rect 53929 11163 53987 11169
rect 54205 11203 54263 11209
rect 54205 11169 54217 11203
rect 54251 11200 54263 11203
rect 54478 11200 54484 11212
rect 54251 11172 54484 11200
rect 54251 11169 54263 11172
rect 54205 11163 54263 11169
rect 54478 11160 54484 11172
rect 54536 11200 54542 11212
rect 54536 11172 55812 11200
rect 54536 11160 54542 11172
rect 51074 11132 51080 11144
rect 50755 11104 51080 11132
rect 50755 11101 50767 11104
rect 50709 11095 50767 11101
rect 47452 11036 47716 11064
rect 47780 11064 47808 11092
rect 49694 11064 49700 11076
rect 47780 11036 49700 11064
rect 47452 11024 47458 11036
rect 49694 11024 49700 11036
rect 49752 11024 49758 11076
rect 50062 11024 50068 11076
rect 50120 11064 50126 11076
rect 50632 11064 50660 11095
rect 51074 11092 51080 11104
rect 51132 11092 51138 11144
rect 51534 11092 51540 11144
rect 51592 11132 51598 11144
rect 51905 11135 51963 11141
rect 51905 11132 51917 11135
rect 51592 11104 51917 11132
rect 51592 11092 51598 11104
rect 51905 11101 51917 11104
rect 51951 11101 51963 11135
rect 51905 11095 51963 11101
rect 51994 11092 52000 11144
rect 52052 11132 52058 11144
rect 52181 11135 52239 11141
rect 52052 11104 52097 11132
rect 52052 11092 52058 11104
rect 52181 11101 52193 11135
rect 52227 11101 52239 11135
rect 52181 11095 52239 11101
rect 52365 11135 52423 11141
rect 52365 11101 52377 11135
rect 52411 11132 52423 11135
rect 53006 11132 53012 11144
rect 52411 11104 53012 11132
rect 52411 11101 52423 11104
rect 52365 11095 52423 11101
rect 50120 11036 50752 11064
rect 50120 11024 50126 11036
rect 50724 11008 50752 11036
rect 51626 11024 51632 11076
rect 51684 11064 51690 11076
rect 52086 11064 52092 11076
rect 51684 11036 52092 11064
rect 51684 11024 51690 11036
rect 52086 11024 52092 11036
rect 52144 11064 52150 11076
rect 52196 11064 52224 11095
rect 53006 11092 53012 11104
rect 53064 11092 53070 11144
rect 53098 11092 53104 11144
rect 53156 11132 53162 11144
rect 54021 11135 54079 11141
rect 54021 11132 54033 11135
rect 53156 11104 54033 11132
rect 53156 11092 53162 11104
rect 54021 11101 54033 11104
rect 54067 11101 54079 11135
rect 54021 11095 54079 11101
rect 52144 11036 52224 11064
rect 53193 11067 53251 11073
rect 52144 11024 52150 11036
rect 53193 11033 53205 11067
rect 53239 11064 53251 11067
rect 53282 11064 53288 11076
rect 53239 11036 53288 11064
rect 53239 11033 53251 11036
rect 53193 11027 53251 11033
rect 53282 11024 53288 11036
rect 53340 11024 53346 11076
rect 54036 11064 54064 11095
rect 54110 11092 54116 11144
rect 54168 11132 54174 11144
rect 54168 11104 54213 11132
rect 54168 11092 54174 11104
rect 55030 11092 55036 11144
rect 55088 11132 55094 11144
rect 55493 11135 55551 11141
rect 55493 11132 55505 11135
rect 55088 11104 55505 11132
rect 55088 11092 55094 11104
rect 55493 11101 55505 11104
rect 55539 11101 55551 11135
rect 55493 11095 55551 11101
rect 54386 11064 54392 11076
rect 54036 11036 54392 11064
rect 54386 11024 54392 11036
rect 54444 11024 54450 11076
rect 54846 11064 54852 11076
rect 54807 11036 54852 11064
rect 54846 11024 54852 11036
rect 54904 11024 54910 11076
rect 43990 10996 43996 11008
rect 43088 10968 43996 10996
rect 43990 10956 43996 10968
rect 44048 10956 44054 11008
rect 44082 10956 44088 11008
rect 44140 10996 44146 11008
rect 45833 10999 45891 11005
rect 45833 10996 45845 10999
rect 44140 10968 45845 10996
rect 44140 10956 44146 10968
rect 45833 10965 45845 10968
rect 45879 10996 45891 10999
rect 45922 10996 45928 11008
rect 45879 10968 45928 10996
rect 45879 10965 45891 10968
rect 45833 10959 45891 10965
rect 45922 10956 45928 10968
rect 45980 10956 45986 11008
rect 47765 10999 47823 11005
rect 47765 10965 47777 10999
rect 47811 10996 47823 10999
rect 48038 10996 48044 11008
rect 47811 10968 48044 10996
rect 47811 10965 47823 10968
rect 47765 10959 47823 10965
rect 48038 10956 48044 10968
rect 48096 10956 48102 11008
rect 48222 10956 48228 11008
rect 48280 10996 48286 11008
rect 50522 10996 50528 11008
rect 48280 10968 50528 10996
rect 48280 10956 48286 10968
rect 50522 10956 50528 10968
rect 50580 10956 50586 11008
rect 50706 10956 50712 11008
rect 50764 10956 50770 11008
rect 50890 10956 50896 11008
rect 50948 10996 50954 11008
rect 52546 10996 52552 11008
rect 50948 10968 52552 10996
rect 50948 10956 50954 10968
rect 52546 10956 52552 10968
rect 52604 10956 52610 11008
rect 52993 10999 53051 11005
rect 52993 10965 53005 10999
rect 53039 10996 53051 10999
rect 53098 10996 53104 11008
rect 53039 10968 53104 10996
rect 53039 10965 53051 10968
rect 52993 10959 53051 10965
rect 53098 10956 53104 10968
rect 53156 10956 53162 11008
rect 53558 10956 53564 11008
rect 53616 10996 53622 11008
rect 55048 10996 55076 11092
rect 55306 11024 55312 11076
rect 55364 11064 55370 11076
rect 55674 11064 55680 11076
rect 55364 11036 55680 11064
rect 55364 11024 55370 11036
rect 55674 11024 55680 11036
rect 55732 11024 55738 11076
rect 55784 11064 55812 11172
rect 55876 11132 55904 11299
rect 58066 11296 58072 11308
rect 58124 11296 58130 11348
rect 56321 11135 56379 11141
rect 56321 11132 56333 11135
rect 55876 11104 56333 11132
rect 56321 11101 56333 11104
rect 56367 11101 56379 11135
rect 56321 11095 56379 11101
rect 56505 11135 56563 11141
rect 56505 11101 56517 11135
rect 56551 11101 56563 11135
rect 56505 11095 56563 11101
rect 56413 11067 56471 11073
rect 56413 11064 56425 11067
rect 55784 11036 56425 11064
rect 56413 11033 56425 11036
rect 56459 11033 56471 11067
rect 56413 11027 56471 11033
rect 56520 11008 56548 11095
rect 53616 10968 55076 10996
rect 53616 10956 53622 10968
rect 55766 10956 55772 11008
rect 55824 10996 55830 11008
rect 56502 10996 56508 11008
rect 55824 10968 56508 10996
rect 55824 10956 55830 10968
rect 56502 10956 56508 10968
rect 56560 10956 56566 11008
rect 56686 10956 56692 11008
rect 56744 10996 56750 11008
rect 56965 10999 57023 11005
rect 56965 10996 56977 10999
rect 56744 10968 56977 10996
rect 56744 10956 56750 10968
rect 56965 10965 56977 10968
rect 57011 10965 57023 10999
rect 57514 10996 57520 11008
rect 57475 10968 57520 10996
rect 56965 10959 57023 10965
rect 57514 10956 57520 10968
rect 57572 10956 57578 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 24486 10752 24492 10804
rect 24544 10792 24550 10804
rect 28721 10795 28779 10801
rect 24544 10764 28212 10792
rect 24544 10752 24550 10764
rect 24213 10727 24271 10733
rect 24213 10693 24225 10727
rect 24259 10724 24271 10727
rect 25222 10724 25228 10736
rect 24259 10696 25228 10724
rect 24259 10693 24271 10696
rect 24213 10687 24271 10693
rect 25222 10684 25228 10696
rect 25280 10684 25286 10736
rect 26418 10724 26424 10736
rect 26252 10696 26424 10724
rect 24762 10616 24768 10668
rect 24820 10656 24826 10668
rect 26252 10665 26280 10696
rect 26418 10684 26424 10696
rect 26476 10724 26482 10736
rect 27430 10724 27436 10736
rect 26476 10696 27436 10724
rect 26476 10684 26482 10696
rect 27430 10684 27436 10696
rect 27488 10684 27494 10736
rect 24949 10659 25007 10665
rect 24949 10656 24961 10659
rect 24820 10628 24961 10656
rect 24820 10616 24826 10628
rect 24949 10625 24961 10628
rect 24995 10625 25007 10659
rect 24949 10619 25007 10625
rect 26237 10659 26295 10665
rect 26237 10625 26249 10659
rect 26283 10625 26295 10659
rect 27338 10656 27344 10668
rect 27299 10628 27344 10656
rect 26237 10619 26295 10625
rect 27338 10616 27344 10628
rect 27396 10616 27402 10668
rect 27614 10656 27620 10668
rect 27575 10628 27620 10656
rect 27614 10616 27620 10628
rect 27672 10616 27678 10668
rect 28184 10656 28212 10764
rect 28721 10761 28733 10795
rect 28767 10792 28779 10795
rect 28767 10764 28994 10792
rect 28767 10761 28779 10764
rect 28721 10755 28779 10761
rect 28626 10724 28632 10736
rect 28587 10696 28632 10724
rect 28626 10684 28632 10696
rect 28684 10684 28690 10736
rect 28966 10724 28994 10764
rect 29454 10752 29460 10804
rect 29512 10792 29518 10804
rect 29914 10792 29920 10804
rect 29512 10764 29920 10792
rect 29512 10752 29518 10764
rect 29914 10752 29920 10764
rect 29972 10752 29978 10804
rect 30282 10792 30288 10804
rect 30243 10764 30288 10792
rect 30282 10752 30288 10764
rect 30340 10752 30346 10804
rect 30374 10752 30380 10804
rect 30432 10792 30438 10804
rect 30742 10792 30748 10804
rect 30432 10764 30748 10792
rect 30432 10752 30438 10764
rect 30742 10752 30748 10764
rect 30800 10752 30806 10804
rect 30926 10752 30932 10804
rect 30984 10792 30990 10804
rect 31021 10795 31079 10801
rect 31021 10792 31033 10795
rect 30984 10764 31033 10792
rect 30984 10752 30990 10764
rect 31021 10761 31033 10764
rect 31067 10761 31079 10795
rect 31021 10755 31079 10761
rect 31294 10752 31300 10804
rect 31352 10792 31358 10804
rect 31352 10764 31432 10792
rect 31352 10752 31358 10764
rect 31404 10733 31432 10764
rect 32030 10752 32036 10804
rect 32088 10792 32094 10804
rect 32309 10795 32367 10801
rect 32309 10792 32321 10795
rect 32088 10764 32321 10792
rect 32088 10752 32094 10764
rect 32309 10761 32321 10764
rect 32355 10761 32367 10795
rect 32309 10755 32367 10761
rect 33686 10752 33692 10804
rect 33744 10792 33750 10804
rect 33873 10795 33931 10801
rect 33873 10792 33885 10795
rect 33744 10764 33885 10792
rect 33744 10752 33750 10764
rect 33873 10761 33885 10764
rect 33919 10761 33931 10795
rect 33873 10755 33931 10761
rect 34606 10752 34612 10804
rect 34664 10792 34670 10804
rect 35069 10795 35127 10801
rect 35069 10792 35081 10795
rect 34664 10764 35081 10792
rect 34664 10752 34670 10764
rect 35069 10761 35081 10764
rect 35115 10761 35127 10795
rect 35069 10755 35127 10761
rect 35342 10752 35348 10804
rect 35400 10792 35406 10804
rect 38197 10795 38255 10801
rect 35400 10764 35572 10792
rect 35400 10752 35406 10764
rect 31189 10727 31247 10733
rect 28966 10696 30236 10724
rect 29178 10656 29184 10668
rect 28184 10628 29184 10656
rect 29178 10616 29184 10628
rect 29236 10616 29242 10668
rect 29825 10659 29883 10665
rect 29825 10625 29837 10659
rect 29871 10625 29883 10659
rect 29825 10619 29883 10625
rect 24670 10588 24676 10600
rect 24631 10560 24676 10588
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 26970 10548 26976 10600
rect 27028 10588 27034 10600
rect 27433 10591 27491 10597
rect 27433 10588 27445 10591
rect 27028 10560 27445 10588
rect 27028 10548 27034 10560
rect 27433 10557 27445 10560
rect 27479 10588 27491 10591
rect 27479 10560 28764 10588
rect 27479 10557 27491 10560
rect 27433 10551 27491 10557
rect 24765 10523 24823 10529
rect 24765 10489 24777 10523
rect 24811 10520 24823 10523
rect 27338 10520 27344 10532
rect 24811 10492 27344 10520
rect 24811 10489 24823 10492
rect 24765 10483 24823 10489
rect 27338 10480 27344 10492
rect 27396 10480 27402 10532
rect 27525 10523 27583 10529
rect 27525 10489 27537 10523
rect 27571 10489 27583 10523
rect 28736 10520 28764 10560
rect 28810 10548 28816 10600
rect 28868 10588 28874 10600
rect 28868 10560 28913 10588
rect 28868 10548 28874 10560
rect 29270 10520 29276 10532
rect 28736 10492 29276 10520
rect 27525 10483 27583 10489
rect 24854 10412 24860 10464
rect 24912 10452 24918 10464
rect 24912 10424 24957 10452
rect 24912 10412 24918 10424
rect 25222 10412 25228 10464
rect 25280 10452 25286 10464
rect 25685 10455 25743 10461
rect 25685 10452 25697 10455
rect 25280 10424 25697 10452
rect 25280 10412 25286 10424
rect 25685 10421 25697 10424
rect 25731 10421 25743 10455
rect 25685 10415 25743 10421
rect 26421 10455 26479 10461
rect 26421 10421 26433 10455
rect 26467 10452 26479 10455
rect 26510 10452 26516 10464
rect 26467 10424 26516 10452
rect 26467 10421 26479 10424
rect 26421 10415 26479 10421
rect 26510 10412 26516 10424
rect 26568 10412 26574 10464
rect 26786 10412 26792 10464
rect 26844 10452 26850 10464
rect 27157 10455 27215 10461
rect 27157 10452 27169 10455
rect 26844 10424 27169 10452
rect 26844 10412 26850 10424
rect 27157 10421 27169 10424
rect 27203 10421 27215 10455
rect 27157 10415 27215 10421
rect 27246 10412 27252 10464
rect 27304 10452 27310 10464
rect 27540 10452 27568 10483
rect 29270 10480 29276 10492
rect 29328 10480 29334 10532
rect 29840 10520 29868 10619
rect 29914 10616 29920 10668
rect 29972 10656 29978 10668
rect 30098 10665 30104 10668
rect 30081 10659 30104 10665
rect 29972 10628 30017 10656
rect 29972 10616 29978 10628
rect 30081 10625 30093 10659
rect 30081 10619 30104 10625
rect 30098 10616 30104 10619
rect 30156 10616 30162 10668
rect 30208 10600 30236 10696
rect 31189 10693 31201 10727
rect 31235 10724 31247 10727
rect 31389 10727 31447 10733
rect 31235 10696 31340 10724
rect 31235 10693 31247 10696
rect 31189 10687 31247 10693
rect 31312 10656 31340 10696
rect 31389 10693 31401 10727
rect 31435 10724 31447 10727
rect 32766 10724 32772 10736
rect 31435 10696 32772 10724
rect 31435 10693 31447 10696
rect 31389 10687 31447 10693
rect 32766 10684 32772 10696
rect 32824 10684 32830 10736
rect 33042 10684 33048 10736
rect 33100 10724 33106 10736
rect 33100 10696 35480 10724
rect 33100 10684 33106 10696
rect 31754 10656 31760 10668
rect 31312 10628 31760 10656
rect 31754 10616 31760 10628
rect 31812 10656 31818 10668
rect 32585 10659 32643 10665
rect 32585 10656 32597 10659
rect 31812 10628 32597 10656
rect 31812 10616 31818 10628
rect 32585 10625 32597 10628
rect 32631 10625 32643 10659
rect 32585 10619 32643 10625
rect 33870 10616 33876 10668
rect 33928 10656 33934 10668
rect 34149 10659 34207 10665
rect 34149 10656 34161 10659
rect 33928 10628 34161 10656
rect 33928 10616 33934 10628
rect 34149 10625 34161 10628
rect 34195 10625 34207 10659
rect 34149 10619 34207 10625
rect 34348 10600 34376 10696
rect 34606 10616 34612 10668
rect 34664 10656 34670 10668
rect 35452 10665 35480 10696
rect 35544 10665 35572 10764
rect 38197 10761 38209 10795
rect 38243 10792 38255 10795
rect 38378 10792 38384 10804
rect 38243 10764 38384 10792
rect 38243 10761 38255 10764
rect 38197 10755 38255 10761
rect 38378 10752 38384 10764
rect 38436 10752 38442 10804
rect 39301 10795 39359 10801
rect 39301 10761 39313 10795
rect 39347 10792 39359 10795
rect 40218 10792 40224 10804
rect 39347 10764 40224 10792
rect 39347 10761 39359 10764
rect 39301 10755 39359 10761
rect 40218 10752 40224 10764
rect 40276 10752 40282 10804
rect 46842 10792 46848 10804
rect 45940 10764 46848 10792
rect 36354 10684 36360 10736
rect 36412 10724 36418 10736
rect 37642 10724 37648 10736
rect 36412 10696 37648 10724
rect 36412 10684 36418 10696
rect 37642 10684 37648 10696
rect 37700 10724 37706 10736
rect 37700 10696 37780 10724
rect 37700 10684 37706 10696
rect 35437 10659 35495 10665
rect 34664 10628 35388 10656
rect 34664 10616 34670 10628
rect 30190 10548 30196 10600
rect 30248 10588 30254 10600
rect 32493 10591 32551 10597
rect 32493 10588 32505 10591
rect 30248 10560 32505 10588
rect 30248 10548 30254 10560
rect 32493 10557 32505 10560
rect 32539 10557 32551 10591
rect 32493 10551 32551 10557
rect 32677 10591 32735 10597
rect 32677 10557 32689 10591
rect 32723 10557 32735 10591
rect 32677 10551 32735 10557
rect 32214 10520 32220 10532
rect 29840 10492 32220 10520
rect 32214 10480 32220 10492
rect 32272 10520 32278 10532
rect 32582 10520 32588 10532
rect 32272 10492 32588 10520
rect 32272 10480 32278 10492
rect 32582 10480 32588 10492
rect 32640 10480 32646 10532
rect 32692 10520 32720 10551
rect 32766 10548 32772 10600
rect 32824 10588 32830 10600
rect 34057 10591 34115 10597
rect 32824 10560 32869 10588
rect 32824 10548 32830 10560
rect 34057 10557 34069 10591
rect 34103 10557 34115 10591
rect 34238 10588 34244 10600
rect 34199 10560 34244 10588
rect 34057 10551 34115 10557
rect 34072 10520 34100 10551
rect 34238 10548 34244 10560
rect 34296 10548 34302 10600
rect 34330 10548 34336 10600
rect 34388 10588 34394 10600
rect 35250 10588 35256 10600
rect 34388 10560 34433 10588
rect 35211 10560 35256 10588
rect 34388 10548 34394 10560
rect 35250 10548 35256 10560
rect 35308 10548 35314 10600
rect 35360 10597 35388 10628
rect 35437 10625 35449 10659
rect 35483 10625 35495 10659
rect 35437 10619 35495 10625
rect 35529 10659 35587 10665
rect 35529 10625 35541 10659
rect 35575 10625 35587 10659
rect 35529 10619 35587 10625
rect 36446 10616 36452 10668
rect 36504 10656 36510 10668
rect 36541 10659 36599 10665
rect 36541 10656 36553 10659
rect 36504 10628 36553 10656
rect 36504 10616 36510 10628
rect 36541 10625 36553 10628
rect 36587 10625 36599 10659
rect 36541 10619 36599 10625
rect 36909 10659 36967 10665
rect 36909 10625 36921 10659
rect 36955 10625 36967 10659
rect 36909 10619 36967 10625
rect 35345 10591 35403 10597
rect 35345 10557 35357 10591
rect 35391 10588 35403 10591
rect 35894 10588 35900 10600
rect 35391 10560 35900 10588
rect 35391 10557 35403 10560
rect 35345 10551 35403 10557
rect 35894 10548 35900 10560
rect 35952 10548 35958 10600
rect 36924 10588 36952 10619
rect 37274 10616 37280 10668
rect 37332 10656 37338 10668
rect 37752 10665 37780 10696
rect 37826 10684 37832 10736
rect 37884 10724 37890 10736
rect 41782 10724 41788 10736
rect 37884 10696 40342 10724
rect 40972 10696 41788 10724
rect 37884 10684 37890 10696
rect 37553 10659 37611 10665
rect 37553 10656 37565 10659
rect 37332 10628 37565 10656
rect 37332 10616 37338 10628
rect 37553 10625 37565 10628
rect 37599 10625 37611 10659
rect 37553 10619 37611 10625
rect 37737 10659 37795 10665
rect 37737 10625 37749 10659
rect 37783 10625 37795 10659
rect 38562 10656 38568 10668
rect 38523 10628 38568 10656
rect 37737 10619 37795 10625
rect 38562 10616 38568 10628
rect 38620 10616 38626 10668
rect 38930 10616 38936 10668
rect 38988 10656 38994 10668
rect 39209 10659 39267 10665
rect 39209 10656 39221 10659
rect 38988 10628 39221 10656
rect 38988 10616 38994 10628
rect 39209 10625 39221 10628
rect 39255 10625 39267 10659
rect 39390 10656 39396 10668
rect 39351 10628 39396 10656
rect 39209 10619 39267 10625
rect 39390 10616 39396 10628
rect 39448 10616 39454 10668
rect 40678 10656 40684 10668
rect 40591 10628 40684 10656
rect 40678 10616 40684 10628
rect 40736 10656 40742 10668
rect 40972 10656 41000 10696
rect 41782 10684 41788 10696
rect 41840 10684 41846 10736
rect 42334 10684 42340 10736
rect 42392 10724 42398 10736
rect 42797 10727 42855 10733
rect 42797 10724 42809 10727
rect 42392 10696 42809 10724
rect 42392 10684 42398 10696
rect 42797 10693 42809 10696
rect 42843 10693 42855 10727
rect 42797 10687 42855 10693
rect 43438 10684 43444 10736
rect 43496 10724 43502 10736
rect 44082 10724 44088 10736
rect 43496 10696 44088 10724
rect 43496 10684 43502 10696
rect 44082 10684 44088 10696
rect 44140 10684 44146 10736
rect 45554 10724 45560 10736
rect 45296 10696 45560 10724
rect 40736 10628 41000 10656
rect 41233 10659 41291 10665
rect 40736 10616 40742 10628
rect 41233 10625 41245 10659
rect 41279 10656 41291 10659
rect 42426 10656 42432 10668
rect 41279 10628 42432 10656
rect 41279 10625 41291 10628
rect 41233 10619 41291 10625
rect 42426 10616 42432 10628
rect 42484 10616 42490 10668
rect 44266 10656 44272 10668
rect 44227 10628 44272 10656
rect 44266 10616 44272 10628
rect 44324 10616 44330 10668
rect 45296 10665 45324 10696
rect 45554 10684 45560 10696
rect 45612 10684 45618 10736
rect 45281 10659 45339 10665
rect 45281 10625 45293 10659
rect 45327 10625 45339 10659
rect 45281 10619 45339 10625
rect 45465 10659 45523 10665
rect 45465 10625 45477 10659
rect 45511 10656 45523 10659
rect 45940 10656 45968 10764
rect 46842 10752 46848 10764
rect 46900 10752 46906 10804
rect 49421 10795 49479 10801
rect 49421 10792 49433 10795
rect 46952 10764 49433 10792
rect 46124 10696 46888 10724
rect 46124 10668 46152 10696
rect 46106 10656 46112 10668
rect 45511 10628 45968 10656
rect 46067 10628 46112 10656
rect 45511 10625 45523 10628
rect 45465 10619 45523 10625
rect 46106 10616 46112 10628
rect 46164 10616 46170 10668
rect 46290 10616 46296 10668
rect 46348 10656 46354 10668
rect 46477 10659 46535 10665
rect 46477 10656 46489 10659
rect 46348 10628 46489 10656
rect 46348 10616 46354 10628
rect 46477 10625 46489 10628
rect 46523 10656 46535 10659
rect 46658 10656 46664 10668
rect 46523 10628 46664 10656
rect 46523 10625 46535 10628
rect 46477 10619 46535 10625
rect 46658 10616 46664 10628
rect 46716 10616 46722 10668
rect 37645 10591 37703 10597
rect 37645 10588 37657 10591
rect 36924 10560 37657 10588
rect 37645 10557 37657 10560
rect 37691 10588 37703 10591
rect 38286 10588 38292 10600
rect 37691 10560 38292 10588
rect 37691 10557 37703 10560
rect 37645 10551 37703 10557
rect 38286 10548 38292 10560
rect 38344 10588 38350 10600
rect 38381 10591 38439 10597
rect 38381 10588 38393 10591
rect 38344 10560 38393 10588
rect 38344 10548 38350 10560
rect 38381 10557 38393 10560
rect 38427 10557 38439 10591
rect 38381 10551 38439 10557
rect 38470 10548 38476 10600
rect 38528 10588 38534 10600
rect 38657 10591 38715 10597
rect 38528 10560 38573 10588
rect 38528 10548 38534 10560
rect 38657 10557 38669 10591
rect 38703 10588 38715 10591
rect 39298 10588 39304 10600
rect 38703 10560 39304 10588
rect 38703 10557 38715 10560
rect 38657 10551 38715 10557
rect 39298 10548 39304 10560
rect 39356 10588 39362 10600
rect 39758 10588 39764 10600
rect 39356 10560 39764 10588
rect 39356 10548 39362 10560
rect 39758 10548 39764 10560
rect 39816 10548 39822 10600
rect 44453 10591 44511 10597
rect 44453 10557 44465 10591
rect 44499 10588 44511 10591
rect 45646 10588 45652 10600
rect 44499 10560 45652 10588
rect 44499 10557 44511 10560
rect 44453 10551 44511 10557
rect 45646 10548 45652 10560
rect 45704 10588 45710 10600
rect 46201 10591 46259 10597
rect 46201 10588 46213 10591
rect 45704 10560 46213 10588
rect 45704 10548 45710 10560
rect 46201 10557 46213 10560
rect 46247 10588 46259 10591
rect 46566 10588 46572 10600
rect 46247 10560 46572 10588
rect 46247 10557 46259 10560
rect 46201 10551 46259 10557
rect 46566 10548 46572 10560
rect 46624 10548 46630 10600
rect 46753 10591 46811 10597
rect 46753 10557 46765 10591
rect 46799 10557 46811 10591
rect 46860 10588 46888 10696
rect 46952 10665 46980 10764
rect 49421 10761 49433 10764
rect 49467 10761 49479 10795
rect 50525 10795 50583 10801
rect 50525 10792 50537 10795
rect 49421 10755 49479 10761
rect 49804 10764 50537 10792
rect 48038 10724 48044 10736
rect 47999 10696 48044 10724
rect 48038 10684 48044 10696
rect 48096 10684 48102 10736
rect 48685 10727 48743 10733
rect 48685 10693 48697 10727
rect 48731 10724 48743 10727
rect 49804 10724 49832 10764
rect 50525 10761 50537 10764
rect 50571 10761 50583 10795
rect 50525 10755 50583 10761
rect 51074 10752 51080 10804
rect 51132 10792 51138 10804
rect 51132 10764 51856 10792
rect 51132 10752 51138 10764
rect 51718 10724 51724 10736
rect 48731 10696 49832 10724
rect 48731 10693 48743 10696
rect 48685 10687 48743 10693
rect 46937 10659 46995 10665
rect 46937 10625 46949 10659
rect 46983 10625 46995 10659
rect 47762 10656 47768 10668
rect 47723 10628 47768 10656
rect 46937 10619 46995 10625
rect 47762 10616 47768 10628
rect 47820 10616 47826 10668
rect 47857 10659 47915 10665
rect 47857 10625 47869 10659
rect 47903 10625 47915 10659
rect 48056 10656 48084 10684
rect 48593 10659 48651 10665
rect 48593 10656 48605 10659
rect 48056 10628 48605 10656
rect 47857 10619 47915 10625
rect 48593 10625 48605 10628
rect 48639 10625 48651 10659
rect 48866 10656 48872 10668
rect 48827 10628 48872 10656
rect 48593 10619 48651 10625
rect 47872 10588 47900 10619
rect 48866 10616 48872 10628
rect 48924 10616 48930 10668
rect 49804 10665 49832 10696
rect 50356 10696 51724 10724
rect 49789 10659 49847 10665
rect 49789 10625 49801 10659
rect 49835 10625 49847 10659
rect 49789 10619 49847 10625
rect 49694 10588 49700 10600
rect 46860 10560 47900 10588
rect 49655 10560 49700 10588
rect 46753 10551 46811 10557
rect 36357 10523 36415 10529
rect 36357 10520 36369 10523
rect 32692 10492 33456 10520
rect 34072 10492 36369 10520
rect 27304 10424 27568 10452
rect 27304 10412 27310 10424
rect 28074 10412 28080 10464
rect 28132 10452 28138 10464
rect 28261 10455 28319 10461
rect 28261 10452 28273 10455
rect 28132 10424 28273 10452
rect 28132 10412 28138 10424
rect 28261 10421 28273 10424
rect 28307 10421 28319 10455
rect 28261 10415 28319 10421
rect 28534 10412 28540 10464
rect 28592 10452 28598 10464
rect 30926 10452 30932 10464
rect 28592 10424 30932 10452
rect 28592 10412 28598 10424
rect 30926 10412 30932 10424
rect 30984 10412 30990 10464
rect 31202 10412 31208 10464
rect 31260 10461 31266 10464
rect 31260 10452 31272 10461
rect 32692 10452 32720 10492
rect 33428 10461 33456 10492
rect 36357 10489 36369 10492
rect 36403 10489 36415 10523
rect 46474 10520 46480 10532
rect 46435 10492 46480 10520
rect 36357 10483 36415 10489
rect 46474 10480 46480 10492
rect 46532 10480 46538 10532
rect 46658 10480 46664 10532
rect 46716 10520 46722 10532
rect 46768 10520 46796 10551
rect 49694 10548 49700 10560
rect 49752 10548 49758 10600
rect 46716 10492 46796 10520
rect 46716 10480 46722 10492
rect 47026 10480 47032 10532
rect 47084 10520 47090 10532
rect 47765 10523 47823 10529
rect 47765 10520 47777 10523
rect 47084 10492 47777 10520
rect 47084 10480 47090 10492
rect 47765 10489 47777 10492
rect 47811 10489 47823 10523
rect 47765 10483 47823 10489
rect 48869 10523 48927 10529
rect 48869 10489 48881 10523
rect 48915 10520 48927 10523
rect 49510 10520 49516 10532
rect 48915 10492 49516 10520
rect 48915 10489 48927 10492
rect 48869 10483 48927 10489
rect 49510 10480 49516 10492
rect 49568 10480 49574 10532
rect 49804 10520 49832 10619
rect 50154 10616 50160 10668
rect 50212 10656 50218 10668
rect 50356 10665 50384 10696
rect 51718 10684 51724 10696
rect 51776 10684 51782 10736
rect 51828 10724 51856 10764
rect 51994 10752 52000 10804
rect 52052 10792 52058 10804
rect 52181 10795 52239 10801
rect 52181 10792 52193 10795
rect 52052 10764 52193 10792
rect 52052 10752 52058 10764
rect 52181 10761 52193 10764
rect 52227 10761 52239 10795
rect 54018 10792 54024 10804
rect 53979 10764 54024 10792
rect 52181 10755 52239 10761
rect 54018 10752 54024 10764
rect 54076 10752 54082 10804
rect 54202 10752 54208 10804
rect 54260 10792 54266 10804
rect 55033 10795 55091 10801
rect 55033 10792 55045 10795
rect 54260 10764 55045 10792
rect 54260 10752 54266 10764
rect 55033 10761 55045 10764
rect 55079 10761 55091 10795
rect 55033 10755 55091 10761
rect 53006 10724 53012 10736
rect 51828 10696 52684 10724
rect 52919 10696 53012 10724
rect 50249 10659 50307 10665
rect 50249 10656 50261 10659
rect 50212 10628 50261 10656
rect 50212 10616 50218 10628
rect 50249 10625 50261 10628
rect 50295 10625 50307 10659
rect 50249 10619 50307 10625
rect 50341 10659 50399 10665
rect 50341 10625 50353 10659
rect 50387 10625 50399 10659
rect 51626 10656 51632 10668
rect 51587 10628 51632 10656
rect 50341 10619 50399 10625
rect 51626 10616 51632 10628
rect 51684 10616 51690 10668
rect 52086 10656 52092 10668
rect 52047 10628 52092 10656
rect 52086 10616 52092 10628
rect 52144 10616 52150 10668
rect 52178 10616 52184 10668
rect 52236 10656 52242 10668
rect 52273 10659 52331 10665
rect 52273 10656 52285 10659
rect 52236 10628 52285 10656
rect 52236 10616 52242 10628
rect 52273 10625 52285 10628
rect 52319 10625 52331 10659
rect 52273 10619 52331 10625
rect 50522 10588 50528 10600
rect 50483 10560 50528 10588
rect 50522 10548 50528 10560
rect 50580 10548 50586 10600
rect 51350 10548 51356 10600
rect 51408 10588 51414 10600
rect 51537 10591 51595 10597
rect 51537 10588 51549 10591
rect 51408 10560 51549 10588
rect 51408 10548 51414 10560
rect 51537 10557 51549 10560
rect 51583 10588 51595 10591
rect 52454 10588 52460 10600
rect 51583 10560 52460 10588
rect 51583 10557 51595 10560
rect 51537 10551 51595 10557
rect 52454 10548 52460 10560
rect 52512 10548 52518 10600
rect 52656 10588 52684 10696
rect 53006 10684 53012 10696
rect 53064 10724 53070 10736
rect 55048 10724 55076 10755
rect 55122 10752 55128 10804
rect 55180 10792 55186 10804
rect 57425 10795 57483 10801
rect 57425 10792 57437 10795
rect 55180 10764 57437 10792
rect 55180 10752 55186 10764
rect 57425 10761 57437 10764
rect 57471 10792 57483 10795
rect 58250 10792 58256 10804
rect 57471 10764 58256 10792
rect 57471 10761 57483 10764
rect 57425 10755 57483 10761
rect 58250 10752 58256 10764
rect 58308 10752 58314 10804
rect 55490 10724 55496 10736
rect 53064 10696 54616 10724
rect 55048 10696 55496 10724
rect 53064 10684 53070 10696
rect 54588 10668 54616 10696
rect 55490 10684 55496 10696
rect 55548 10724 55554 10736
rect 56318 10724 56324 10736
rect 55548 10696 56324 10724
rect 55548 10684 55554 10696
rect 56318 10684 56324 10696
rect 56376 10684 56382 10736
rect 52914 10656 52920 10668
rect 52875 10628 52920 10656
rect 52914 10616 52920 10628
rect 52972 10616 52978 10668
rect 53101 10659 53159 10665
rect 53101 10625 53113 10659
rect 53147 10656 53159 10659
rect 53282 10656 53288 10668
rect 53147 10628 53288 10656
rect 53147 10625 53159 10628
rect 53101 10619 53159 10625
rect 53116 10588 53144 10619
rect 53282 10616 53288 10628
rect 53340 10616 53346 10668
rect 54202 10656 54208 10668
rect 54163 10628 54208 10656
rect 54202 10616 54208 10628
rect 54260 10616 54266 10668
rect 54294 10616 54300 10668
rect 54352 10656 54358 10668
rect 54570 10656 54576 10668
rect 54352 10628 54397 10656
rect 54531 10628 54576 10656
rect 54352 10616 54358 10628
rect 54570 10616 54576 10628
rect 54628 10616 54634 10668
rect 56134 10616 56140 10668
rect 56192 10656 56198 10668
rect 56229 10659 56287 10665
rect 56229 10656 56241 10659
rect 56192 10628 56241 10656
rect 56192 10616 56198 10628
rect 56229 10625 56241 10628
rect 56275 10625 56287 10659
rect 56229 10619 56287 10625
rect 52656 10560 53144 10588
rect 54312 10520 54340 10616
rect 54478 10588 54484 10600
rect 54439 10560 54484 10588
rect 54478 10548 54484 10560
rect 54536 10548 54542 10600
rect 55953 10523 56011 10529
rect 55953 10520 55965 10523
rect 49804 10492 51488 10520
rect 54312 10492 55965 10520
rect 31260 10424 32720 10452
rect 33413 10455 33471 10461
rect 31260 10415 31272 10424
rect 33413 10421 33425 10455
rect 33459 10452 33471 10455
rect 35526 10452 35532 10464
rect 33459 10424 35532 10452
rect 33459 10421 33471 10424
rect 33413 10415 33471 10421
rect 31260 10412 31266 10415
rect 35526 10412 35532 10424
rect 35584 10412 35590 10464
rect 36722 10452 36728 10464
rect 36683 10424 36728 10452
rect 36722 10412 36728 10424
rect 36780 10412 36786 10464
rect 43070 10412 43076 10464
rect 43128 10452 43134 10464
rect 43257 10455 43315 10461
rect 43257 10452 43269 10455
rect 43128 10424 43269 10452
rect 43128 10412 43134 10424
rect 43257 10421 43269 10424
rect 43303 10452 43315 10455
rect 43714 10452 43720 10464
rect 43303 10424 43720 10452
rect 43303 10421 43315 10424
rect 43257 10415 43315 10421
rect 43714 10412 43720 10424
rect 43772 10412 43778 10464
rect 44082 10452 44088 10464
rect 44043 10424 44088 10452
rect 44082 10412 44088 10424
rect 44140 10412 44146 10464
rect 45370 10452 45376 10464
rect 45331 10424 45376 10452
rect 45370 10412 45376 10424
rect 45428 10412 45434 10464
rect 45830 10412 45836 10464
rect 45888 10452 45894 10464
rect 46934 10452 46940 10464
rect 45888 10424 46940 10452
rect 45888 10412 45894 10424
rect 46934 10412 46940 10424
rect 46992 10452 46998 10464
rect 49418 10452 49424 10464
rect 46992 10424 49424 10452
rect 46992 10412 46998 10424
rect 49418 10412 49424 10424
rect 49476 10412 49482 10464
rect 49786 10452 49792 10464
rect 49747 10424 49792 10452
rect 49786 10412 49792 10424
rect 49844 10412 49850 10464
rect 51261 10455 51319 10461
rect 51261 10421 51273 10455
rect 51307 10452 51319 10455
rect 51350 10452 51356 10464
rect 51307 10424 51356 10452
rect 51307 10421 51319 10424
rect 51261 10415 51319 10421
rect 51350 10412 51356 10424
rect 51408 10412 51414 10464
rect 51460 10461 51488 10492
rect 55953 10489 55965 10492
rect 55999 10489 56011 10523
rect 55953 10483 56011 10489
rect 51445 10455 51503 10461
rect 51445 10421 51457 10455
rect 51491 10421 51503 10455
rect 51445 10415 51503 10421
rect 52638 10412 52644 10464
rect 52696 10452 52702 10464
rect 55306 10452 55312 10464
rect 52696 10424 55312 10452
rect 52696 10412 52702 10424
rect 55306 10412 55312 10424
rect 55364 10412 55370 10464
rect 56778 10452 56784 10464
rect 56739 10424 56784 10452
rect 56778 10412 56784 10424
rect 56836 10412 56842 10464
rect 57974 10412 57980 10464
rect 58032 10452 58038 10464
rect 58069 10455 58127 10461
rect 58069 10452 58081 10455
rect 58032 10424 58081 10452
rect 58032 10412 58038 10424
rect 58069 10421 58081 10424
rect 58115 10421 58127 10455
rect 58069 10415 58127 10421
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 24581 10251 24639 10257
rect 24581 10217 24593 10251
rect 24627 10248 24639 10251
rect 24670 10248 24676 10260
rect 24627 10220 24676 10248
rect 24627 10217 24639 10220
rect 24581 10211 24639 10217
rect 24670 10208 24676 10220
rect 24728 10208 24734 10260
rect 26237 10251 26295 10257
rect 26237 10217 26249 10251
rect 26283 10248 26295 10251
rect 26326 10248 26332 10260
rect 26283 10220 26332 10248
rect 26283 10217 26295 10220
rect 26237 10211 26295 10217
rect 26326 10208 26332 10220
rect 26384 10208 26390 10260
rect 26786 10248 26792 10260
rect 26747 10220 26792 10248
rect 26786 10208 26792 10220
rect 26844 10208 26850 10260
rect 27706 10208 27712 10260
rect 27764 10248 27770 10260
rect 27982 10248 27988 10260
rect 27764 10220 27988 10248
rect 27764 10208 27770 10220
rect 27982 10208 27988 10220
rect 28040 10208 28046 10260
rect 28442 10248 28448 10260
rect 28403 10220 28448 10248
rect 28442 10208 28448 10220
rect 28500 10208 28506 10260
rect 28626 10208 28632 10260
rect 28684 10248 28690 10260
rect 28902 10248 28908 10260
rect 28684 10220 28908 10248
rect 28684 10208 28690 10220
rect 28902 10208 28908 10220
rect 28960 10208 28966 10260
rect 29178 10248 29184 10260
rect 29139 10220 29184 10248
rect 29178 10208 29184 10220
rect 29236 10248 29242 10260
rect 29822 10248 29828 10260
rect 29236 10220 29828 10248
rect 29236 10208 29242 10220
rect 29822 10208 29828 10220
rect 29880 10208 29886 10260
rect 29917 10251 29975 10257
rect 29917 10217 29929 10251
rect 29963 10248 29975 10251
rect 30190 10248 30196 10260
rect 29963 10220 30196 10248
rect 29963 10217 29975 10220
rect 29917 10211 29975 10217
rect 30190 10208 30196 10220
rect 30248 10208 30254 10260
rect 30558 10248 30564 10260
rect 30519 10220 30564 10248
rect 30558 10208 30564 10220
rect 30616 10208 30622 10260
rect 31573 10251 31631 10257
rect 31573 10217 31585 10251
rect 31619 10248 31631 10251
rect 31754 10248 31760 10260
rect 31619 10220 31760 10248
rect 31619 10217 31631 10220
rect 31573 10211 31631 10217
rect 31754 10208 31760 10220
rect 31812 10208 31818 10260
rect 33134 10208 33140 10260
rect 33192 10248 33198 10260
rect 33778 10248 33784 10260
rect 33192 10220 33784 10248
rect 33192 10208 33198 10220
rect 33778 10208 33784 10220
rect 33836 10248 33842 10260
rect 36446 10248 36452 10260
rect 33836 10220 36452 10248
rect 33836 10208 33842 10220
rect 36446 10208 36452 10220
rect 36504 10208 36510 10260
rect 37550 10208 37556 10260
rect 37608 10248 37614 10260
rect 38289 10251 38347 10257
rect 38289 10248 38301 10251
rect 37608 10220 38301 10248
rect 37608 10208 37614 10220
rect 38289 10217 38301 10220
rect 38335 10217 38347 10251
rect 38289 10211 38347 10217
rect 38473 10251 38531 10257
rect 38473 10217 38485 10251
rect 38519 10248 38531 10251
rect 38654 10248 38660 10260
rect 38519 10220 38660 10248
rect 38519 10217 38531 10220
rect 38473 10211 38531 10217
rect 38654 10208 38660 10220
rect 38712 10208 38718 10260
rect 38746 10208 38752 10260
rect 38804 10248 38810 10260
rect 38933 10251 38991 10257
rect 38933 10248 38945 10251
rect 38804 10220 38945 10248
rect 38804 10208 38810 10220
rect 38933 10217 38945 10220
rect 38979 10217 38991 10251
rect 43165 10251 43223 10257
rect 43165 10248 43177 10251
rect 38933 10211 38991 10217
rect 42260 10220 43177 10248
rect 28534 10140 28540 10192
rect 28592 10180 28598 10192
rect 28592 10152 34284 10180
rect 28592 10140 28598 10152
rect 25222 10112 25228 10124
rect 24044 10084 25228 10112
rect 23842 10044 23848 10056
rect 23803 10016 23848 10044
rect 23842 10004 23848 10016
rect 23900 10004 23906 10056
rect 24044 10053 24072 10084
rect 25222 10072 25228 10084
rect 25280 10072 25286 10124
rect 27154 10072 27160 10124
rect 27212 10112 27218 10124
rect 32493 10115 32551 10121
rect 27212 10084 28258 10112
rect 27212 10072 27218 10084
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10013 24087 10047
rect 24854 10044 24860 10056
rect 24815 10016 24860 10044
rect 24029 10007 24087 10013
rect 24854 10004 24860 10016
rect 24912 10044 24918 10056
rect 25317 10047 25375 10053
rect 25317 10044 25329 10047
rect 24912 10016 25329 10044
rect 24912 10004 24918 10016
rect 25317 10013 25329 10016
rect 25363 10013 25375 10047
rect 25317 10007 25375 10013
rect 25501 10047 25559 10053
rect 25501 10013 25513 10047
rect 25547 10013 25559 10047
rect 25501 10007 25559 10013
rect 25777 10047 25835 10053
rect 25777 10013 25789 10047
rect 25823 10044 25835 10047
rect 25958 10044 25964 10056
rect 25823 10016 25964 10044
rect 25823 10013 25835 10016
rect 25777 10007 25835 10013
rect 24578 9976 24584 9988
rect 24539 9948 24584 9976
rect 24578 9936 24584 9948
rect 24636 9936 24642 9988
rect 24762 9976 24768 9988
rect 24723 9948 24768 9976
rect 24762 9936 24768 9948
rect 24820 9936 24826 9988
rect 25516 9976 25544 10007
rect 25958 10004 25964 10016
rect 26016 10004 26022 10056
rect 26418 10047 26476 10053
rect 26418 10013 26430 10047
rect 26464 10044 26476 10047
rect 26602 10044 26608 10056
rect 26464 10016 26608 10044
rect 26464 10013 26476 10016
rect 26418 10007 26476 10013
rect 26602 10004 26608 10016
rect 26660 10004 26666 10056
rect 26878 10044 26884 10056
rect 26839 10016 26884 10044
rect 26878 10004 26884 10016
rect 26936 10004 26942 10056
rect 27338 10004 27344 10056
rect 27396 10044 27402 10056
rect 27801 10047 27859 10053
rect 27801 10044 27813 10047
rect 27396 10016 27813 10044
rect 27396 10004 27402 10016
rect 27801 10013 27813 10016
rect 27847 10013 27859 10047
rect 27801 10007 27859 10013
rect 27985 10047 28043 10053
rect 27985 10013 27997 10047
rect 28031 10013 28043 10047
rect 27985 10007 28043 10013
rect 26326 9976 26332 9988
rect 25516 9948 26332 9976
rect 26326 9936 26332 9948
rect 26384 9936 26390 9988
rect 28000 9976 28028 10007
rect 28074 10004 28080 10056
rect 28132 10044 28138 10056
rect 28230 10053 28258 10084
rect 30392 10084 31432 10112
rect 28215 10047 28273 10053
rect 28132 10016 28177 10044
rect 28132 10004 28138 10016
rect 28215 10013 28227 10047
rect 28261 10044 28273 10047
rect 28810 10044 28816 10056
rect 28261 10016 28816 10044
rect 28261 10013 28273 10016
rect 28215 10007 28273 10013
rect 28810 10004 28816 10016
rect 28868 10004 28874 10056
rect 29086 10004 29092 10056
rect 29144 10044 29150 10056
rect 29733 10047 29791 10053
rect 29733 10044 29745 10047
rect 29144 10016 29745 10044
rect 29144 10004 29150 10016
rect 29733 10013 29745 10016
rect 29779 10013 29791 10047
rect 29733 10007 29791 10013
rect 29822 10004 29828 10056
rect 29880 10044 29886 10056
rect 29917 10047 29975 10053
rect 29917 10044 29929 10047
rect 29880 10016 29929 10044
rect 29880 10004 29886 10016
rect 29917 10013 29929 10016
rect 29963 10044 29975 10047
rect 30098 10044 30104 10056
rect 29963 10016 30104 10044
rect 29963 10013 29975 10016
rect 29917 10007 29975 10013
rect 30098 10004 30104 10016
rect 30156 10004 30162 10056
rect 30392 10053 30420 10084
rect 30377 10047 30435 10053
rect 30377 10013 30389 10047
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 30558 10004 30564 10056
rect 30616 10044 30622 10056
rect 31294 10044 31300 10056
rect 30616 10016 31300 10044
rect 30616 10004 30622 10016
rect 31294 10004 31300 10016
rect 31352 10004 31358 10056
rect 31404 10044 31432 10084
rect 32493 10081 32505 10115
rect 32539 10112 32551 10115
rect 32766 10112 32772 10124
rect 32539 10084 32772 10112
rect 32539 10081 32551 10084
rect 32493 10075 32551 10081
rect 32766 10072 32772 10084
rect 32824 10112 32830 10124
rect 33870 10112 33876 10124
rect 32824 10084 33088 10112
rect 33831 10084 33876 10112
rect 32824 10072 32830 10084
rect 31481 10047 31539 10053
rect 31481 10044 31493 10047
rect 31404 10016 31493 10044
rect 31481 10013 31493 10016
rect 31527 10013 31539 10047
rect 31662 10044 31668 10056
rect 31623 10016 31668 10044
rect 31481 10007 31539 10013
rect 31202 9976 31208 9988
rect 28000 9948 31208 9976
rect 31202 9936 31208 9948
rect 31260 9936 31266 9988
rect 31496 9976 31524 10007
rect 31662 10004 31668 10016
rect 31720 10004 31726 10056
rect 32214 10004 32220 10056
rect 32272 10044 32278 10056
rect 33060 10053 33088 10084
rect 33870 10072 33876 10084
rect 33928 10072 33934 10124
rect 33962 10072 33968 10124
rect 34020 10112 34026 10124
rect 34020 10084 34192 10112
rect 34020 10072 34026 10084
rect 32401 10047 32459 10053
rect 32401 10044 32413 10047
rect 32272 10016 32413 10044
rect 32272 10004 32278 10016
rect 32401 10013 32413 10016
rect 32447 10013 32459 10047
rect 32401 10007 32459 10013
rect 32585 10047 32643 10053
rect 32585 10013 32597 10047
rect 32631 10044 32643 10047
rect 33045 10047 33103 10053
rect 32631 10038 32904 10044
rect 32631 10016 32996 10038
rect 32631 10013 32643 10016
rect 32585 10007 32643 10013
rect 32876 10010 32996 10016
rect 31938 9976 31944 9988
rect 31496 9948 31944 9976
rect 31938 9936 31944 9948
rect 31996 9936 32002 9988
rect 24029 9911 24087 9917
rect 24029 9877 24041 9911
rect 24075 9908 24087 9911
rect 24780 9908 24808 9936
rect 25682 9908 25688 9920
rect 24075 9880 24808 9908
rect 25643 9880 25688 9908
rect 24075 9877 24087 9880
rect 24029 9871 24087 9877
rect 25682 9868 25688 9880
rect 25740 9868 25746 9920
rect 26421 9911 26479 9917
rect 26421 9877 26433 9911
rect 26467 9908 26479 9911
rect 28350 9908 28356 9920
rect 26467 9880 28356 9908
rect 26467 9877 26479 9880
rect 26421 9871 26479 9877
rect 28350 9868 28356 9880
rect 28408 9868 28414 9920
rect 29546 9868 29552 9920
rect 29604 9908 29610 9920
rect 29914 9908 29920 9920
rect 29604 9880 29920 9908
rect 29604 9868 29610 9880
rect 29914 9868 29920 9880
rect 29972 9868 29978 9920
rect 30098 9868 30104 9920
rect 30156 9908 30162 9920
rect 31294 9908 31300 9920
rect 30156 9880 31300 9908
rect 30156 9868 30162 9880
rect 31294 9868 31300 9880
rect 31352 9868 31358 9920
rect 31662 9868 31668 9920
rect 31720 9908 31726 9920
rect 32766 9908 32772 9920
rect 31720 9880 32772 9908
rect 31720 9868 31726 9880
rect 32766 9868 32772 9880
rect 32824 9868 32830 9920
rect 32968 9908 32996 10010
rect 33045 10013 33057 10047
rect 33091 10013 33103 10047
rect 33045 10007 33103 10013
rect 33226 10004 33232 10056
rect 33284 10053 33290 10056
rect 33284 10047 33299 10053
rect 33287 10013 33299 10047
rect 33284 10007 33299 10013
rect 33781 10047 33839 10053
rect 33781 10013 33793 10047
rect 33827 10013 33839 10047
rect 34054 10044 34060 10056
rect 34015 10016 34060 10044
rect 33781 10007 33839 10013
rect 33284 10004 33290 10007
rect 33137 9979 33195 9985
rect 33137 9945 33149 9979
rect 33183 9976 33195 9979
rect 33502 9976 33508 9988
rect 33183 9948 33508 9976
rect 33183 9945 33195 9948
rect 33137 9939 33195 9945
rect 33502 9936 33508 9948
rect 33560 9936 33566 9988
rect 33686 9976 33692 9988
rect 33647 9948 33692 9976
rect 33686 9936 33692 9948
rect 33744 9936 33750 9988
rect 33796 9976 33824 10007
rect 34054 10004 34060 10016
rect 34112 10004 34118 10056
rect 34164 10053 34192 10084
rect 34149 10047 34207 10053
rect 34149 10013 34161 10047
rect 34195 10013 34207 10047
rect 34256 10044 34284 10152
rect 35986 10140 35992 10192
rect 36044 10180 36050 10192
rect 36817 10183 36875 10189
rect 36817 10180 36829 10183
rect 36044 10152 36829 10180
rect 36044 10140 36050 10152
rect 36817 10149 36829 10152
rect 36863 10149 36875 10183
rect 36817 10143 36875 10149
rect 41601 10183 41659 10189
rect 41601 10149 41613 10183
rect 41647 10180 41659 10183
rect 41647 10152 42196 10180
rect 41647 10149 41659 10152
rect 41601 10143 41659 10149
rect 34330 10072 34336 10124
rect 34388 10112 34394 10124
rect 36538 10112 36544 10124
rect 34388 10084 36400 10112
rect 36499 10084 36544 10112
rect 34388 10072 34394 10084
rect 35345 10047 35403 10053
rect 35345 10044 35357 10047
rect 34256 10016 35357 10044
rect 34149 10007 34207 10013
rect 35345 10013 35357 10016
rect 35391 10013 35403 10047
rect 35802 10044 35808 10056
rect 35763 10016 35808 10044
rect 35345 10007 35403 10013
rect 35802 10004 35808 10016
rect 35860 10004 35866 10056
rect 36372 10053 36400 10084
rect 36538 10072 36544 10084
rect 36596 10072 36602 10124
rect 41230 10112 41236 10124
rect 40236 10084 41236 10112
rect 40236 10056 40264 10084
rect 41230 10072 41236 10084
rect 41288 10072 41294 10124
rect 42168 10121 42196 10152
rect 42153 10115 42211 10121
rect 42153 10081 42165 10115
rect 42199 10081 42211 10115
rect 42153 10075 42211 10081
rect 36357 10047 36415 10053
rect 36357 10013 36369 10047
rect 36403 10044 36415 10047
rect 36906 10044 36912 10056
rect 36403 10016 36492 10044
rect 36867 10016 36912 10044
rect 36403 10013 36415 10016
rect 36357 10007 36415 10013
rect 36170 9976 36176 9988
rect 33796 9948 36176 9976
rect 36170 9936 36176 9948
rect 36228 9936 36234 9988
rect 34330 9908 34336 9920
rect 32968 9880 34336 9908
rect 34330 9868 34336 9880
rect 34388 9908 34394 9920
rect 34606 9908 34612 9920
rect 34388 9880 34612 9908
rect 34388 9868 34394 9880
rect 34606 9868 34612 9880
rect 34664 9868 34670 9920
rect 34790 9868 34796 9920
rect 34848 9908 34854 9920
rect 35802 9908 35808 9920
rect 34848 9880 35808 9908
rect 34848 9868 34854 9880
rect 35802 9868 35808 9880
rect 35860 9868 35866 9920
rect 36464 9908 36492 10016
rect 36906 10004 36912 10016
rect 36964 10004 36970 10056
rect 38838 10004 38844 10056
rect 38896 10044 38902 10056
rect 39114 10044 39120 10056
rect 38896 10016 39120 10044
rect 38896 10004 38902 10016
rect 39114 10004 39120 10016
rect 39172 10004 39178 10056
rect 39206 10004 39212 10056
rect 39264 10044 39270 10056
rect 40037 10047 40095 10053
rect 40037 10044 40049 10047
rect 39264 10016 40049 10044
rect 39264 10004 39270 10016
rect 40037 10013 40049 10016
rect 40083 10013 40095 10047
rect 40218 10044 40224 10056
rect 40179 10016 40224 10044
rect 40037 10007 40095 10013
rect 40218 10004 40224 10016
rect 40276 10004 40282 10056
rect 41322 10044 41328 10056
rect 41283 10016 41328 10044
rect 41322 10004 41328 10016
rect 41380 10004 41386 10056
rect 42260 10053 42288 10220
rect 43165 10217 43177 10220
rect 43211 10248 43223 10251
rect 43809 10251 43867 10257
rect 43809 10248 43821 10251
rect 43211 10220 43821 10248
rect 43211 10217 43223 10220
rect 43165 10211 43223 10217
rect 43809 10217 43821 10220
rect 43855 10217 43867 10251
rect 43809 10211 43867 10217
rect 43993 10251 44051 10257
rect 43993 10217 44005 10251
rect 44039 10248 44051 10251
rect 45646 10248 45652 10260
rect 44039 10220 45652 10248
rect 44039 10217 44051 10220
rect 43993 10211 44051 10217
rect 45646 10208 45652 10220
rect 45704 10208 45710 10260
rect 45922 10248 45928 10260
rect 45883 10220 45928 10248
rect 45922 10208 45928 10220
rect 45980 10208 45986 10260
rect 46106 10208 46112 10260
rect 46164 10248 46170 10260
rect 47213 10251 47271 10257
rect 47213 10248 47225 10251
rect 46164 10220 47225 10248
rect 46164 10208 46170 10220
rect 47213 10217 47225 10220
rect 47259 10217 47271 10251
rect 47670 10248 47676 10260
rect 47631 10220 47676 10248
rect 47213 10211 47271 10217
rect 47670 10208 47676 10220
rect 47728 10208 47734 10260
rect 49145 10251 49203 10257
rect 49145 10217 49157 10251
rect 49191 10248 49203 10251
rect 49234 10248 49240 10260
rect 49191 10220 49240 10248
rect 49191 10217 49203 10220
rect 49145 10211 49203 10217
rect 49234 10208 49240 10220
rect 49292 10208 49298 10260
rect 49418 10208 49424 10260
rect 49476 10248 49482 10260
rect 50430 10248 50436 10260
rect 49476 10220 50436 10248
rect 49476 10208 49482 10220
rect 50430 10208 50436 10220
rect 50488 10208 50494 10260
rect 50801 10251 50859 10257
rect 50801 10217 50813 10251
rect 50847 10248 50859 10251
rect 51626 10248 51632 10260
rect 50847 10220 51632 10248
rect 50847 10217 50859 10220
rect 50801 10211 50859 10217
rect 51626 10208 51632 10220
rect 51684 10208 51690 10260
rect 52178 10208 52184 10260
rect 52236 10248 52242 10260
rect 52365 10251 52423 10257
rect 52365 10248 52377 10251
rect 52236 10220 52377 10248
rect 52236 10208 52242 10220
rect 52365 10217 52377 10220
rect 52411 10248 52423 10251
rect 52638 10248 52644 10260
rect 52411 10220 52644 10248
rect 52411 10217 52423 10220
rect 52365 10211 52423 10217
rect 52638 10208 52644 10220
rect 52696 10208 52702 10260
rect 53098 10208 53104 10260
rect 53156 10248 53162 10260
rect 53193 10251 53251 10257
rect 53193 10248 53205 10251
rect 53156 10220 53205 10248
rect 53156 10208 53162 10220
rect 53193 10217 53205 10220
rect 53239 10248 53251 10251
rect 53742 10248 53748 10260
rect 53239 10220 53748 10248
rect 53239 10217 53251 10220
rect 53193 10211 53251 10217
rect 53742 10208 53748 10220
rect 53800 10208 53806 10260
rect 53837 10251 53895 10257
rect 53837 10217 53849 10251
rect 53883 10248 53895 10251
rect 54110 10248 54116 10260
rect 53883 10220 54116 10248
rect 53883 10217 53895 10220
rect 53837 10211 53895 10217
rect 54110 10208 54116 10220
rect 54168 10208 54174 10260
rect 54481 10251 54539 10257
rect 54481 10217 54493 10251
rect 54527 10248 54539 10251
rect 56686 10248 56692 10260
rect 54527 10220 56692 10248
rect 54527 10217 54539 10220
rect 54481 10211 54539 10217
rect 42613 10183 42671 10189
rect 42613 10149 42625 10183
rect 42659 10180 42671 10183
rect 42659 10152 45324 10180
rect 42659 10149 42671 10152
rect 42613 10143 42671 10149
rect 45296 10121 45324 10152
rect 45370 10140 45376 10192
rect 45428 10180 45434 10192
rect 47949 10183 48007 10189
rect 47949 10180 47961 10183
rect 45428 10152 47961 10180
rect 45428 10140 45434 10152
rect 47949 10149 47961 10152
rect 47995 10180 48007 10183
rect 48866 10180 48872 10192
rect 47995 10152 48872 10180
rect 47995 10149 48007 10152
rect 47949 10143 48007 10149
rect 48866 10140 48872 10152
rect 48924 10140 48930 10192
rect 50154 10180 50160 10192
rect 49344 10152 50160 10180
rect 43349 10115 43407 10121
rect 43349 10081 43361 10115
rect 43395 10112 43407 10115
rect 45281 10115 45339 10121
rect 43395 10084 45232 10112
rect 43395 10081 43407 10084
rect 43349 10075 43407 10081
rect 42245 10047 42303 10053
rect 42245 10013 42257 10047
rect 42291 10013 42303 10047
rect 42245 10007 42303 10013
rect 43073 10047 43131 10053
rect 43073 10013 43085 10047
rect 43119 10044 43131 10047
rect 44082 10044 44088 10056
rect 43119 10016 44088 10044
rect 43119 10013 43131 10016
rect 43073 10007 43131 10013
rect 44082 10004 44088 10016
rect 44140 10004 44146 10056
rect 44358 10004 44364 10056
rect 44416 10004 44422 10056
rect 36538 9936 36544 9988
rect 36596 9976 36602 9988
rect 36998 9976 37004 9988
rect 36596 9948 37004 9976
rect 36596 9936 36602 9948
rect 36998 9936 37004 9948
rect 37056 9936 37062 9988
rect 38102 9976 38108 9988
rect 38063 9948 38108 9976
rect 38102 9936 38108 9948
rect 38160 9936 38166 9988
rect 38286 9936 38292 9988
rect 38344 9985 38350 9988
rect 38344 9979 38363 9985
rect 38351 9945 38363 9979
rect 40402 9976 40408 9988
rect 40363 9948 40408 9976
rect 38344 9939 38363 9945
rect 38344 9936 38350 9939
rect 40402 9936 40408 9948
rect 40460 9936 40466 9988
rect 41601 9979 41659 9985
rect 41601 9945 41613 9979
rect 41647 9976 41659 9979
rect 43162 9976 43168 9988
rect 41647 9948 43168 9976
rect 41647 9945 41659 9948
rect 41601 9939 41659 9945
rect 43162 9936 43168 9948
rect 43220 9936 43226 9988
rect 43346 9976 43352 9988
rect 43307 9948 43352 9976
rect 43346 9936 43352 9948
rect 43404 9936 43410 9988
rect 43990 9985 43996 9988
rect 43977 9979 43996 9985
rect 43977 9945 43989 9979
rect 43977 9939 43996 9945
rect 43990 9936 43996 9939
rect 44048 9936 44054 9988
rect 44177 9979 44235 9985
rect 44177 9945 44189 9979
rect 44223 9976 44235 9979
rect 44376 9976 44404 10004
rect 44542 9976 44548 9988
rect 44223 9948 44548 9976
rect 44223 9945 44235 9948
rect 44177 9939 44235 9945
rect 44542 9936 44548 9948
rect 44600 9936 44606 9988
rect 45204 9976 45232 10084
rect 45281 10081 45293 10115
rect 45327 10081 45339 10115
rect 45281 10075 45339 10081
rect 46750 10072 46756 10124
rect 46808 10112 46814 10124
rect 48041 10115 48099 10121
rect 46808 10084 47900 10112
rect 46808 10072 46814 10084
rect 45738 10044 45744 10056
rect 45702 10016 45744 10044
rect 45738 10004 45744 10016
rect 45796 10004 45802 10056
rect 46842 10044 46848 10056
rect 46803 10016 46848 10044
rect 46842 10004 46848 10016
rect 46900 10004 46906 10056
rect 47872 10053 47900 10084
rect 48041 10081 48053 10115
rect 48087 10112 48099 10115
rect 48682 10112 48688 10124
rect 48087 10084 48688 10112
rect 48087 10081 48099 10084
rect 48041 10075 48099 10081
rect 48682 10072 48688 10084
rect 48740 10072 48746 10124
rect 49344 10121 49372 10152
rect 50154 10140 50160 10152
rect 50212 10140 50218 10192
rect 50448 10180 50476 10208
rect 50890 10180 50896 10192
rect 50448 10152 50896 10180
rect 50890 10140 50896 10152
rect 50948 10140 50954 10192
rect 51442 10180 51448 10192
rect 51403 10152 51448 10180
rect 51442 10140 51448 10152
rect 51500 10140 51506 10192
rect 51534 10140 51540 10192
rect 51592 10180 51598 10192
rect 51592 10152 51637 10180
rect 51592 10140 51598 10152
rect 51718 10140 51724 10192
rect 51776 10180 51782 10192
rect 51994 10180 52000 10192
rect 51776 10152 52000 10180
rect 51776 10140 51782 10152
rect 51994 10140 52000 10152
rect 52052 10180 52058 10192
rect 52052 10152 53144 10180
rect 52052 10140 52058 10152
rect 49329 10115 49387 10121
rect 49329 10081 49341 10115
rect 49375 10081 49387 10115
rect 53006 10112 53012 10124
rect 49329 10075 49387 10081
rect 49712 10084 53012 10112
rect 47029 10047 47087 10053
rect 47029 10013 47041 10047
rect 47075 10013 47087 10047
rect 47029 10007 47087 10013
rect 47857 10047 47915 10053
rect 47857 10013 47869 10047
rect 47903 10013 47915 10047
rect 48130 10044 48136 10056
rect 48091 10016 48136 10044
rect 47857 10007 47915 10013
rect 45922 9976 45928 9988
rect 45204 9948 45928 9976
rect 45922 9936 45928 9948
rect 45980 9936 45986 9988
rect 46198 9936 46204 9988
rect 46256 9976 46262 9988
rect 46750 9976 46756 9988
rect 46256 9948 46756 9976
rect 46256 9936 46262 9948
rect 46750 9936 46756 9948
rect 46808 9936 46814 9988
rect 40420 9908 40448 9936
rect 36464 9880 40448 9908
rect 41417 9911 41475 9917
rect 41417 9877 41429 9911
rect 41463 9908 41475 9911
rect 43438 9908 43444 9920
rect 41463 9880 43444 9908
rect 41463 9877 41475 9880
rect 41417 9871 41475 9877
rect 43438 9868 43444 9880
rect 43496 9868 43502 9920
rect 45738 9908 45744 9920
rect 45699 9880 45744 9908
rect 45738 9868 45744 9880
rect 45796 9868 45802 9920
rect 47044 9908 47072 10007
rect 47872 9976 47900 10007
rect 48130 10004 48136 10016
rect 48188 10004 48194 10056
rect 48317 10047 48375 10053
rect 48317 10013 48329 10047
rect 48363 10044 48375 10047
rect 49050 10044 49056 10056
rect 48363 10016 49056 10044
rect 48363 10013 48375 10016
rect 48317 10007 48375 10013
rect 49050 10004 49056 10016
rect 49108 10004 49114 10056
rect 49418 10044 49424 10056
rect 49379 10016 49424 10044
rect 49418 10004 49424 10016
rect 49476 10004 49482 10056
rect 49712 9985 49740 10084
rect 53006 10072 53012 10084
rect 53064 10072 53070 10124
rect 53116 10112 53144 10152
rect 53282 10140 53288 10192
rect 53340 10180 53346 10192
rect 54496 10180 54524 10211
rect 56686 10208 56692 10220
rect 56744 10208 56750 10260
rect 53340 10152 54524 10180
rect 53340 10140 53346 10152
rect 55674 10140 55680 10192
rect 55732 10180 55738 10192
rect 58161 10183 58219 10189
rect 58161 10180 58173 10183
rect 55732 10152 58173 10180
rect 55732 10140 55738 10152
rect 58161 10149 58173 10152
rect 58207 10149 58219 10183
rect 58161 10143 58219 10149
rect 56778 10112 56784 10124
rect 53116 10084 56784 10112
rect 50430 10004 50436 10056
rect 50488 10044 50494 10056
rect 50617 10047 50675 10053
rect 50617 10044 50629 10047
rect 50488 10016 50629 10044
rect 50488 10004 50494 10016
rect 50617 10013 50629 10016
rect 50663 10013 50675 10047
rect 50798 10044 50804 10056
rect 50759 10016 50804 10044
rect 50617 10007 50675 10013
rect 50798 10004 50804 10016
rect 50856 10004 50862 10056
rect 51350 10044 51356 10056
rect 51311 10016 51356 10044
rect 51350 10004 51356 10016
rect 51408 10004 51414 10056
rect 51626 10044 51632 10056
rect 51587 10016 51632 10044
rect 51626 10004 51632 10016
rect 51684 10004 51690 10056
rect 53098 10044 53104 10056
rect 53059 10016 53104 10044
rect 53098 10004 53104 10016
rect 53156 10004 53162 10056
rect 53300 10053 53328 10084
rect 56778 10072 56784 10084
rect 56836 10072 56842 10124
rect 53285 10047 53343 10053
rect 53285 10013 53297 10047
rect 53331 10013 53343 10047
rect 53285 10007 53343 10013
rect 53742 10004 53748 10056
rect 53800 10044 53806 10056
rect 53929 10047 53987 10053
rect 53800 10016 53845 10044
rect 53800 10004 53806 10016
rect 53929 10013 53941 10047
rect 53975 10013 53987 10047
rect 56134 10044 56140 10056
rect 56095 10016 56140 10044
rect 53929 10007 53987 10013
rect 49697 9979 49755 9985
rect 49697 9976 49709 9979
rect 47872 9948 49709 9976
rect 49697 9945 49709 9948
rect 49743 9945 49755 9979
rect 49697 9939 49755 9945
rect 49786 9936 49792 9988
rect 49844 9976 49850 9988
rect 50816 9976 50844 10004
rect 49844 9948 50844 9976
rect 51813 9979 51871 9985
rect 49844 9936 49850 9948
rect 51813 9945 51825 9979
rect 51859 9976 51871 9979
rect 53834 9976 53840 9988
rect 51859 9948 53840 9976
rect 51859 9945 51871 9948
rect 51813 9939 51871 9945
rect 53834 9936 53840 9948
rect 53892 9936 53898 9988
rect 50706 9908 50712 9920
rect 47044 9880 50712 9908
rect 50706 9868 50712 9880
rect 50764 9868 50770 9920
rect 53098 9868 53104 9920
rect 53156 9908 53162 9920
rect 53466 9908 53472 9920
rect 53156 9880 53472 9908
rect 53156 9868 53162 9880
rect 53466 9868 53472 9880
rect 53524 9868 53530 9920
rect 53742 9868 53748 9920
rect 53800 9908 53806 9920
rect 53944 9908 53972 10007
rect 56134 10004 56140 10016
rect 56192 10004 56198 10056
rect 56410 10044 56416 10056
rect 56371 10016 56416 10044
rect 56410 10004 56416 10016
rect 56468 10004 56474 10056
rect 57238 10004 57244 10056
rect 57296 10044 57302 10056
rect 57974 10044 57980 10056
rect 57296 10016 57980 10044
rect 57296 10004 57302 10016
rect 57974 10004 57980 10016
rect 58032 10004 58038 10056
rect 57422 9976 57428 9988
rect 55968 9948 57428 9976
rect 53800 9880 53972 9908
rect 53800 9868 53806 9880
rect 55306 9868 55312 9920
rect 55364 9908 55370 9920
rect 55968 9917 55996 9948
rect 57422 9936 57428 9948
rect 57480 9936 57486 9988
rect 55953 9911 56011 9917
rect 55953 9908 55965 9911
rect 55364 9880 55965 9908
rect 55364 9868 55370 9880
rect 55953 9877 55965 9880
rect 55999 9877 56011 9911
rect 55953 9871 56011 9877
rect 56962 9868 56968 9920
rect 57020 9908 57026 9920
rect 57057 9911 57115 9917
rect 57057 9908 57069 9911
rect 57020 9880 57069 9908
rect 57020 9868 57026 9880
rect 57057 9877 57069 9880
rect 57103 9877 57115 9911
rect 57057 9871 57115 9877
rect 57146 9868 57152 9920
rect 57204 9908 57210 9920
rect 57606 9908 57612 9920
rect 57204 9880 57612 9908
rect 57204 9868 57210 9880
rect 57606 9868 57612 9880
rect 57664 9868 57670 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 26878 9664 26884 9716
rect 26936 9704 26942 9716
rect 27433 9707 27491 9713
rect 27433 9704 27445 9707
rect 26936 9676 27445 9704
rect 26936 9664 26942 9676
rect 27433 9673 27445 9676
rect 27479 9673 27491 9707
rect 27433 9667 27491 9673
rect 28810 9664 28816 9716
rect 28868 9704 28874 9716
rect 28868 9676 31340 9704
rect 28868 9664 28874 9676
rect 23753 9639 23811 9645
rect 23753 9605 23765 9639
rect 23799 9636 23811 9639
rect 24118 9636 24124 9648
rect 23799 9608 24124 9636
rect 23799 9605 23811 9608
rect 23753 9599 23811 9605
rect 24118 9596 24124 9608
rect 24176 9636 24182 9648
rect 24857 9639 24915 9645
rect 24857 9636 24869 9639
rect 24176 9608 24869 9636
rect 24176 9596 24182 9608
rect 24857 9605 24869 9608
rect 24903 9636 24915 9639
rect 25774 9636 25780 9648
rect 24903 9608 25780 9636
rect 24903 9605 24915 9608
rect 24857 9599 24915 9605
rect 25774 9596 25780 9608
rect 25832 9596 25838 9648
rect 26786 9596 26792 9648
rect 26844 9636 26850 9648
rect 27246 9636 27252 9648
rect 26844 9608 27252 9636
rect 26844 9596 26850 9608
rect 27246 9596 27252 9608
rect 27304 9596 27310 9648
rect 27341 9639 27399 9645
rect 27341 9605 27353 9639
rect 27387 9636 27399 9639
rect 27798 9636 27804 9648
rect 27387 9608 27804 9636
rect 27387 9605 27399 9608
rect 27341 9599 27399 9605
rect 27798 9596 27804 9608
rect 27856 9596 27862 9648
rect 28350 9596 28356 9648
rect 28408 9636 28414 9648
rect 28445 9639 28503 9645
rect 28445 9636 28457 9639
rect 28408 9608 28457 9636
rect 28408 9596 28414 9608
rect 28445 9605 28457 9608
rect 28491 9605 28503 9639
rect 28445 9599 28503 9605
rect 28534 9596 28540 9648
rect 28592 9636 28598 9648
rect 30745 9639 30803 9645
rect 28592 9608 28764 9636
rect 28592 9596 28598 9608
rect 25958 9528 25964 9580
rect 26016 9568 26022 9580
rect 27890 9568 27896 9580
rect 26016 9540 27896 9568
rect 26016 9528 26022 9540
rect 27890 9528 27896 9540
rect 27948 9528 27954 9580
rect 28258 9528 28264 9580
rect 28316 9528 28322 9580
rect 28626 9568 28632 9580
rect 28587 9540 28632 9568
rect 28626 9528 28632 9540
rect 28684 9528 28690 9580
rect 28736 9577 28764 9608
rect 29472 9608 30236 9636
rect 28721 9571 28779 9577
rect 28721 9537 28733 9571
rect 28767 9537 28779 9571
rect 28721 9531 28779 9537
rect 28905 9571 28963 9577
rect 28905 9537 28917 9571
rect 28951 9537 28963 9571
rect 29472 9568 29500 9608
rect 28905 9531 28963 9537
rect 29007 9561 29065 9567
rect 24305 9503 24363 9509
rect 24305 9469 24317 9503
rect 24351 9500 24363 9503
rect 24578 9500 24584 9512
rect 24351 9472 24584 9500
rect 24351 9469 24363 9472
rect 24305 9463 24363 9469
rect 24578 9460 24584 9472
rect 24636 9500 24642 9512
rect 26053 9503 26111 9509
rect 26053 9500 26065 9503
rect 24636 9472 26065 9500
rect 24636 9460 24642 9472
rect 26053 9469 26065 9472
rect 26099 9500 26111 9503
rect 26602 9500 26608 9512
rect 26099 9472 26608 9500
rect 26099 9469 26111 9472
rect 26053 9463 26111 9469
rect 26602 9460 26608 9472
rect 26660 9500 26666 9512
rect 27614 9500 27620 9512
rect 26660 9472 27620 9500
rect 26660 9460 26666 9472
rect 27614 9460 27620 9472
rect 27672 9460 27678 9512
rect 27709 9503 27767 9509
rect 27709 9469 27721 9503
rect 27755 9500 27767 9503
rect 28276 9500 28304 9528
rect 27755 9472 28304 9500
rect 27755 9469 27767 9472
rect 27709 9463 27767 9469
rect 28810 9460 28816 9512
rect 28868 9500 28874 9512
rect 28920 9500 28948 9531
rect 29007 9527 29019 9561
rect 29053 9558 29065 9561
rect 29196 9558 29500 9568
rect 29053 9540 29500 9558
rect 29053 9530 29224 9540
rect 29053 9527 29065 9530
rect 29546 9528 29552 9580
rect 29604 9568 29610 9580
rect 29641 9571 29699 9577
rect 29641 9568 29653 9571
rect 29604 9540 29653 9568
rect 29604 9528 29610 9540
rect 29641 9537 29653 9540
rect 29687 9537 29699 9571
rect 29822 9568 29828 9580
rect 29783 9540 29828 9568
rect 29641 9531 29699 9537
rect 29822 9528 29828 9540
rect 29880 9528 29886 9580
rect 30098 9568 30104 9580
rect 30059 9540 30104 9568
rect 30098 9528 30104 9540
rect 30156 9528 30162 9580
rect 30208 9568 30236 9608
rect 30745 9605 30757 9639
rect 30791 9636 30803 9639
rect 31110 9636 31116 9648
rect 30791 9608 31116 9636
rect 30791 9605 30803 9608
rect 30745 9599 30803 9605
rect 31110 9596 31116 9608
rect 31168 9596 31174 9648
rect 30926 9568 30932 9580
rect 30208 9540 30932 9568
rect 30926 9528 30932 9540
rect 30984 9528 30990 9580
rect 31021 9571 31079 9577
rect 31021 9537 31033 9571
rect 31067 9537 31079 9571
rect 31202 9568 31208 9580
rect 31163 9540 31208 9568
rect 31021 9531 31079 9537
rect 29007 9521 29065 9527
rect 28868 9472 28948 9500
rect 29917 9503 29975 9509
rect 28868 9460 28874 9472
rect 29917 9469 29929 9503
rect 29963 9500 29975 9503
rect 30006 9500 30012 9512
rect 29963 9472 30012 9500
rect 29963 9469 29975 9472
rect 29917 9463 29975 9469
rect 30006 9460 30012 9472
rect 30064 9500 30070 9512
rect 30558 9500 30564 9512
rect 30064 9472 30564 9500
rect 30064 9460 30070 9472
rect 30558 9460 30564 9472
rect 30616 9460 30622 9512
rect 31036 9500 31064 9531
rect 31202 9528 31208 9540
rect 31260 9528 31266 9580
rect 31312 9577 31340 9676
rect 33870 9664 33876 9716
rect 33928 9704 33934 9716
rect 34149 9707 34207 9713
rect 34149 9704 34161 9707
rect 33928 9676 34161 9704
rect 33928 9664 33934 9676
rect 34149 9673 34161 9676
rect 34195 9673 34207 9707
rect 36357 9707 36415 9713
rect 34149 9667 34207 9673
rect 34992 9676 36308 9704
rect 31570 9596 31576 9648
rect 31628 9636 31634 9648
rect 32398 9636 32404 9648
rect 31628 9608 32404 9636
rect 31628 9596 31634 9608
rect 32398 9596 32404 9608
rect 32456 9596 32462 9648
rect 32674 9596 32680 9648
rect 32732 9636 32738 9648
rect 32769 9639 32827 9645
rect 32769 9636 32781 9639
rect 32732 9608 32781 9636
rect 32732 9596 32738 9608
rect 32769 9605 32781 9608
rect 32815 9605 32827 9639
rect 32769 9599 32827 9605
rect 32950 9577 32956 9614
rect 31297 9571 31355 9577
rect 31297 9537 31309 9571
rect 31343 9537 31355 9571
rect 31297 9531 31355 9537
rect 32936 9571 32956 9577
rect 32936 9537 32948 9571
rect 33008 9562 33014 9614
rect 34054 9596 34060 9648
rect 34112 9636 34118 9648
rect 34992 9636 35020 9676
rect 34112 9608 35020 9636
rect 35989 9639 36047 9645
rect 34112 9596 34118 9608
rect 32982 9540 32996 9562
rect 32982 9537 32994 9540
rect 32936 9531 32994 9537
rect 33042 9528 33048 9580
rect 33100 9568 33106 9580
rect 33318 9568 33324 9580
rect 33100 9540 33145 9568
rect 33279 9540 33324 9568
rect 33100 9528 33106 9540
rect 33318 9528 33324 9540
rect 33376 9528 33382 9580
rect 33781 9571 33839 9577
rect 33781 9537 33793 9571
rect 33827 9568 33839 9571
rect 33870 9568 33876 9580
rect 33827 9540 33876 9568
rect 33827 9537 33839 9540
rect 33781 9531 33839 9537
rect 33870 9528 33876 9540
rect 33928 9528 33934 9580
rect 34900 9577 34928 9608
rect 35989 9605 36001 9639
rect 36035 9636 36047 9639
rect 36035 9608 36069 9636
rect 36035 9605 36047 9608
rect 35989 9599 36047 9605
rect 33965 9571 34023 9577
rect 33965 9537 33977 9571
rect 34011 9568 34023 9571
rect 34885 9571 34943 9577
rect 34011 9540 34192 9568
rect 34011 9537 34023 9540
rect 33965 9531 34023 9537
rect 32030 9500 32036 9512
rect 31036 9472 32036 9500
rect 32030 9460 32036 9472
rect 32088 9460 32094 9512
rect 27525 9435 27583 9441
rect 27525 9401 27537 9435
rect 27571 9432 27583 9435
rect 29362 9432 29368 9444
rect 27571 9404 29368 9432
rect 27571 9401 27583 9404
rect 27525 9395 27583 9401
rect 29362 9392 29368 9404
rect 29420 9392 29426 9444
rect 29457 9435 29515 9441
rect 29457 9401 29469 9435
rect 29503 9432 29515 9435
rect 29638 9432 29644 9444
rect 29503 9404 29644 9432
rect 29503 9401 29515 9404
rect 29457 9395 29515 9401
rect 29638 9392 29644 9404
rect 29696 9392 29702 9444
rect 29733 9435 29791 9441
rect 29733 9401 29745 9435
rect 29779 9401 29791 9435
rect 29733 9395 29791 9401
rect 24946 9364 24952 9376
rect 24907 9336 24952 9364
rect 24946 9324 24952 9336
rect 25004 9364 25010 9376
rect 26418 9364 26424 9376
rect 25004 9336 26424 9364
rect 25004 9324 25010 9336
rect 26418 9324 26424 9336
rect 26476 9324 26482 9376
rect 26605 9367 26663 9373
rect 26605 9333 26617 9367
rect 26651 9364 26663 9367
rect 27246 9364 27252 9376
rect 26651 9336 27252 9364
rect 26651 9333 26663 9336
rect 26605 9327 26663 9333
rect 27246 9324 27252 9336
rect 27304 9324 27310 9376
rect 27617 9367 27675 9373
rect 27617 9333 27629 9367
rect 27663 9364 27675 9367
rect 27706 9364 27712 9376
rect 27663 9336 27712 9364
rect 27663 9333 27675 9336
rect 27617 9327 27675 9333
rect 27706 9324 27712 9336
rect 27764 9324 27770 9376
rect 28350 9324 28356 9376
rect 28408 9364 28414 9376
rect 29748 9364 29776 9395
rect 30098 9392 30104 9444
rect 30156 9432 30162 9444
rect 30650 9432 30656 9444
rect 30156 9404 30656 9432
rect 30156 9392 30162 9404
rect 30650 9392 30656 9404
rect 30708 9392 30714 9444
rect 31110 9392 31116 9444
rect 31168 9432 31174 9444
rect 33134 9432 33140 9444
rect 31168 9404 33140 9432
rect 31168 9392 31174 9404
rect 33134 9392 33140 9404
rect 33192 9392 33198 9444
rect 33229 9435 33287 9441
rect 33229 9401 33241 9435
rect 33275 9432 33287 9435
rect 33502 9432 33508 9444
rect 33275 9404 33508 9432
rect 33275 9401 33287 9404
rect 33229 9395 33287 9401
rect 33502 9392 33508 9404
rect 33560 9392 33566 9444
rect 28408 9336 29776 9364
rect 28408 9324 28414 9336
rect 31294 9324 31300 9376
rect 31352 9364 31358 9376
rect 34054 9364 34060 9376
rect 31352 9336 34060 9364
rect 31352 9324 31358 9336
rect 34054 9324 34060 9336
rect 34112 9324 34118 9376
rect 34164 9364 34192 9540
rect 34885 9537 34897 9571
rect 34931 9568 34943 9571
rect 35069 9571 35127 9577
rect 34931 9540 34965 9568
rect 34931 9537 34943 9540
rect 34885 9531 34943 9537
rect 35069 9537 35081 9571
rect 35115 9568 35127 9571
rect 36004 9568 36032 9599
rect 36170 9596 36176 9648
rect 36228 9645 36234 9648
rect 36228 9639 36247 9645
rect 36235 9605 36247 9639
rect 36280 9636 36308 9676
rect 36357 9673 36369 9707
rect 36403 9704 36415 9707
rect 36906 9704 36912 9716
rect 36403 9676 36912 9704
rect 36403 9673 36415 9676
rect 36357 9667 36415 9673
rect 36906 9664 36912 9676
rect 36964 9664 36970 9716
rect 39758 9704 39764 9716
rect 37476 9676 37872 9704
rect 39719 9676 39764 9704
rect 36280 9608 36676 9636
rect 36228 9599 36247 9605
rect 36228 9596 36234 9599
rect 36538 9568 36544 9580
rect 35115 9540 36544 9568
rect 35115 9537 35127 9540
rect 35069 9531 35127 9537
rect 36538 9528 36544 9540
rect 36596 9528 36602 9580
rect 36648 9568 36676 9608
rect 37274 9568 37280 9580
rect 36648 9540 37280 9568
rect 37274 9528 37280 9540
rect 37332 9528 37338 9580
rect 37476 9577 37504 9676
rect 37844 9636 37872 9676
rect 39758 9664 39764 9676
rect 39816 9664 39822 9716
rect 44266 9664 44272 9716
rect 44324 9704 44330 9716
rect 45462 9704 45468 9716
rect 44324 9676 45468 9704
rect 44324 9664 44330 9676
rect 45462 9664 45468 9676
rect 45520 9704 45526 9716
rect 46474 9704 46480 9716
rect 45520 9676 46480 9704
rect 45520 9664 45526 9676
rect 46474 9664 46480 9676
rect 46532 9664 46538 9716
rect 48590 9664 48596 9716
rect 48648 9704 48654 9716
rect 49326 9704 49332 9716
rect 48648 9676 49332 9704
rect 48648 9664 48654 9676
rect 49326 9664 49332 9676
rect 49384 9704 49390 9716
rect 52086 9704 52092 9716
rect 49384 9676 52092 9704
rect 49384 9664 49390 9676
rect 52086 9664 52092 9676
rect 52144 9664 52150 9716
rect 56134 9664 56140 9716
rect 56192 9704 56198 9716
rect 56321 9707 56379 9713
rect 56321 9704 56333 9707
rect 56192 9676 56333 9704
rect 56192 9664 56198 9676
rect 56321 9673 56333 9676
rect 56367 9673 56379 9707
rect 56321 9667 56379 9673
rect 56410 9664 56416 9716
rect 56468 9664 56474 9716
rect 39390 9636 39396 9648
rect 37844 9608 39396 9636
rect 39390 9596 39396 9608
rect 39448 9636 39454 9648
rect 40865 9639 40923 9645
rect 40865 9636 40877 9639
rect 39448 9608 40877 9636
rect 39448 9596 39454 9608
rect 40865 9605 40877 9608
rect 40911 9605 40923 9639
rect 44358 9636 44364 9648
rect 44319 9608 44364 9636
rect 40865 9599 40923 9605
rect 44358 9596 44364 9608
rect 44416 9596 44422 9648
rect 44545 9639 44603 9645
rect 44545 9605 44557 9639
rect 44591 9636 44603 9639
rect 45649 9639 45707 9645
rect 45649 9636 45661 9639
rect 44591 9608 45661 9636
rect 44591 9605 44603 9608
rect 44545 9599 44603 9605
rect 45649 9605 45661 9608
rect 45695 9605 45707 9639
rect 45649 9599 45707 9605
rect 45922 9596 45928 9648
rect 45980 9636 45986 9648
rect 47118 9636 47124 9648
rect 45980 9608 47124 9636
rect 45980 9596 45986 9608
rect 47118 9596 47124 9608
rect 47176 9596 47182 9648
rect 48682 9636 48688 9648
rect 48643 9608 48688 9636
rect 48682 9596 48688 9608
rect 48740 9596 48746 9648
rect 49234 9636 49240 9648
rect 49160 9608 49240 9636
rect 37461 9571 37519 9577
rect 37461 9537 37473 9571
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 35434 9460 35440 9512
rect 35492 9500 35498 9512
rect 36817 9503 36875 9509
rect 36817 9500 36829 9503
rect 35492 9472 36829 9500
rect 35492 9460 35498 9472
rect 36817 9469 36829 9472
rect 36863 9469 36875 9503
rect 36817 9463 36875 9469
rect 36998 9460 37004 9512
rect 37056 9500 37062 9512
rect 37476 9500 37504 9531
rect 38102 9528 38108 9580
rect 38160 9568 38166 9580
rect 38197 9571 38255 9577
rect 38197 9568 38209 9571
rect 38160 9540 38209 9568
rect 38160 9528 38166 9540
rect 38197 9537 38209 9540
rect 38243 9537 38255 9571
rect 39574 9568 39580 9580
rect 39535 9540 39580 9568
rect 38197 9531 38255 9537
rect 39574 9528 39580 9540
rect 39632 9568 39638 9580
rect 40218 9568 40224 9580
rect 39632 9540 40224 9568
rect 39632 9528 39638 9540
rect 40218 9528 40224 9540
rect 40276 9528 40282 9580
rect 41230 9528 41236 9580
rect 41288 9568 41294 9580
rect 43625 9571 43683 9577
rect 41288 9540 41414 9568
rect 41288 9528 41294 9540
rect 37056 9472 37504 9500
rect 37737 9503 37795 9509
rect 37056 9460 37062 9472
rect 37737 9469 37749 9503
rect 37783 9500 37795 9503
rect 38746 9500 38752 9512
rect 37783 9472 38752 9500
rect 37783 9469 37795 9472
rect 37737 9463 37795 9469
rect 38746 9460 38752 9472
rect 38804 9460 38810 9512
rect 34422 9392 34428 9444
rect 34480 9432 34486 9444
rect 38102 9432 38108 9444
rect 34480 9404 38108 9432
rect 34480 9392 34486 9404
rect 38102 9392 38108 9404
rect 38160 9392 38166 9444
rect 38194 9392 38200 9444
rect 38252 9432 38258 9444
rect 38933 9435 38991 9441
rect 38933 9432 38945 9435
rect 38252 9404 38945 9432
rect 38252 9392 38258 9404
rect 38933 9401 38945 9404
rect 38979 9432 38991 9435
rect 40313 9435 40371 9441
rect 40313 9432 40325 9435
rect 38979 9404 40325 9432
rect 38979 9401 38991 9404
rect 38933 9395 38991 9401
rect 40313 9401 40325 9404
rect 40359 9432 40371 9435
rect 40954 9432 40960 9444
rect 40359 9404 40960 9432
rect 40359 9401 40371 9404
rect 40313 9395 40371 9401
rect 40954 9392 40960 9404
rect 41012 9392 41018 9444
rect 41386 9432 41414 9540
rect 43625 9537 43637 9571
rect 43671 9568 43683 9571
rect 43990 9568 43996 9580
rect 43671 9540 43996 9568
rect 43671 9537 43683 9540
rect 43625 9531 43683 9537
rect 43990 9528 43996 9540
rect 44048 9528 44054 9580
rect 44085 9571 44143 9577
rect 44085 9537 44097 9571
rect 44131 9568 44143 9571
rect 44726 9568 44732 9580
rect 44131 9540 44732 9568
rect 44131 9537 44143 9540
rect 44085 9531 44143 9537
rect 44726 9528 44732 9540
rect 44784 9528 44790 9580
rect 45097 9571 45155 9577
rect 45097 9537 45109 9571
rect 45143 9568 45155 9571
rect 45278 9568 45284 9580
rect 45143 9540 45284 9568
rect 45143 9537 45155 9540
rect 45097 9531 45155 9537
rect 45278 9528 45284 9540
rect 45336 9528 45342 9580
rect 45830 9568 45836 9580
rect 45791 9540 45836 9568
rect 45830 9528 45836 9540
rect 45888 9528 45894 9580
rect 46014 9568 46020 9580
rect 45975 9540 46020 9568
rect 46014 9528 46020 9540
rect 46072 9528 46078 9580
rect 46109 9571 46167 9577
rect 46109 9537 46121 9571
rect 46155 9568 46167 9571
rect 46155 9540 46796 9568
rect 46155 9537 46167 9540
rect 46109 9531 46167 9537
rect 43533 9503 43591 9509
rect 43533 9469 43545 9503
rect 43579 9500 43591 9503
rect 45554 9500 45560 9512
rect 43579 9472 45560 9500
rect 43579 9469 43591 9472
rect 43533 9463 43591 9469
rect 45554 9460 45560 9472
rect 45612 9460 45618 9512
rect 45741 9503 45799 9509
rect 45741 9469 45753 9503
rect 45787 9500 45799 9503
rect 46198 9500 46204 9512
rect 45787 9472 46204 9500
rect 45787 9469 45799 9472
rect 45741 9463 45799 9469
rect 46198 9460 46204 9472
rect 46256 9460 46262 9512
rect 46768 9500 46796 9540
rect 46842 9528 46848 9580
rect 46900 9568 46906 9580
rect 48133 9571 48191 9577
rect 48133 9568 48145 9571
rect 46900 9540 48145 9568
rect 46900 9528 46906 9540
rect 48133 9537 48145 9540
rect 48179 9537 48191 9571
rect 48133 9531 48191 9537
rect 48866 9528 48872 9580
rect 48924 9577 48930 9580
rect 49160 9577 49188 9608
rect 49234 9596 49240 9608
rect 49292 9596 49298 9648
rect 50246 9636 50252 9648
rect 50159 9608 50252 9636
rect 50246 9596 50252 9608
rect 50304 9636 50310 9648
rect 50890 9636 50896 9648
rect 50304 9608 50896 9636
rect 50304 9596 50310 9608
rect 50890 9596 50896 9608
rect 50948 9596 50954 9648
rect 51902 9636 51908 9648
rect 51863 9608 51908 9636
rect 51902 9596 51908 9608
rect 51960 9596 51966 9648
rect 52730 9636 52736 9648
rect 52196 9608 52736 9636
rect 48924 9571 48957 9577
rect 48945 9537 48957 9571
rect 48924 9531 48957 9537
rect 49145 9571 49203 9577
rect 49145 9537 49157 9571
rect 49191 9537 49203 9571
rect 49786 9568 49792 9580
rect 49145 9531 49203 9537
rect 49436 9540 49792 9568
rect 48924 9528 48930 9531
rect 48314 9500 48320 9512
rect 46768 9472 48320 9500
rect 48314 9460 48320 9472
rect 48372 9460 48378 9512
rect 49436 9500 49464 9540
rect 49786 9528 49792 9540
rect 49844 9528 49850 9580
rect 50062 9528 50068 9580
rect 50120 9568 50126 9580
rect 52089 9571 52147 9577
rect 52089 9568 52101 9571
rect 50120 9540 52101 9568
rect 50120 9528 50126 9540
rect 52089 9537 52101 9540
rect 52135 9537 52147 9571
rect 52089 9531 52147 9537
rect 49344 9472 49464 9500
rect 41509 9435 41567 9441
rect 41509 9432 41521 9435
rect 41386 9404 41521 9432
rect 41509 9401 41521 9404
rect 41555 9432 41567 9435
rect 41969 9435 42027 9441
rect 41969 9432 41981 9435
rect 41555 9404 41981 9432
rect 41555 9401 41567 9404
rect 41509 9395 41567 9401
rect 41969 9401 41981 9404
rect 42015 9401 42027 9435
rect 41969 9395 42027 9401
rect 43257 9435 43315 9441
rect 43257 9401 43269 9435
rect 43303 9432 43315 9435
rect 43303 9404 43852 9432
rect 43303 9401 43315 9404
rect 43257 9395 43315 9401
rect 34606 9364 34612 9376
rect 34164 9336 34612 9364
rect 34606 9324 34612 9336
rect 34664 9364 34670 9376
rect 34885 9367 34943 9373
rect 34885 9364 34897 9367
rect 34664 9336 34897 9364
rect 34664 9324 34670 9336
rect 34885 9333 34897 9336
rect 34931 9333 34943 9367
rect 34885 9327 34943 9333
rect 35253 9367 35311 9373
rect 35253 9333 35265 9367
rect 35299 9364 35311 9367
rect 35342 9364 35348 9376
rect 35299 9336 35348 9364
rect 35299 9333 35311 9336
rect 35253 9327 35311 9333
rect 35342 9324 35348 9336
rect 35400 9324 35406 9376
rect 36170 9364 36176 9376
rect 36131 9336 36176 9364
rect 36170 9324 36176 9336
rect 36228 9324 36234 9376
rect 36906 9324 36912 9376
rect 36964 9364 36970 9376
rect 37553 9367 37611 9373
rect 37553 9364 37565 9367
rect 36964 9336 37565 9364
rect 36964 9324 36970 9336
rect 37553 9333 37565 9336
rect 37599 9333 37611 9367
rect 37553 9327 37611 9333
rect 37642 9324 37648 9376
rect 37700 9364 37706 9376
rect 38381 9367 38439 9373
rect 37700 9336 37745 9364
rect 37700 9324 37706 9336
rect 38381 9333 38393 9367
rect 38427 9364 38439 9367
rect 38562 9364 38568 9376
rect 38427 9336 38568 9364
rect 38427 9333 38439 9336
rect 38381 9327 38439 9333
rect 38562 9324 38568 9336
rect 38620 9324 38626 9376
rect 42426 9324 42432 9376
rect 42484 9364 42490 9376
rect 42610 9364 42616 9376
rect 42484 9336 42616 9364
rect 42484 9324 42490 9336
rect 42610 9324 42616 9336
rect 42668 9324 42674 9376
rect 43625 9367 43683 9373
rect 43625 9333 43637 9367
rect 43671 9364 43683 9367
rect 43714 9364 43720 9376
rect 43671 9336 43720 9364
rect 43671 9333 43683 9336
rect 43625 9327 43683 9333
rect 43714 9324 43720 9336
rect 43772 9324 43778 9376
rect 43824 9364 43852 9404
rect 46474 9392 46480 9444
rect 46532 9432 46538 9444
rect 47949 9435 48007 9441
rect 46532 9404 47256 9432
rect 46532 9392 46538 9404
rect 44334 9367 44392 9373
rect 44334 9364 44346 9367
rect 43824 9336 44346 9364
rect 44334 9333 44346 9336
rect 44380 9333 44392 9367
rect 44334 9327 44392 9333
rect 46661 9367 46719 9373
rect 46661 9333 46673 9367
rect 46707 9364 46719 9367
rect 46934 9364 46940 9376
rect 46707 9336 46940 9364
rect 46707 9333 46719 9336
rect 46661 9327 46719 9333
rect 46934 9324 46940 9336
rect 46992 9324 46998 9376
rect 47228 9373 47256 9404
rect 47949 9401 47961 9435
rect 47995 9432 48007 9435
rect 48130 9432 48136 9444
rect 47995 9404 48136 9432
rect 47995 9401 48007 9404
rect 47949 9395 48007 9401
rect 48130 9392 48136 9404
rect 48188 9432 48194 9444
rect 48958 9432 48964 9444
rect 48188 9404 48964 9432
rect 48188 9392 48194 9404
rect 48958 9392 48964 9404
rect 49016 9392 49022 9444
rect 49053 9435 49111 9441
rect 49053 9401 49065 9435
rect 49099 9432 49111 9435
rect 49344 9432 49372 9472
rect 49099 9404 49372 9432
rect 49697 9435 49755 9441
rect 49099 9401 49111 9404
rect 49053 9395 49111 9401
rect 49697 9401 49709 9435
rect 49743 9432 49755 9435
rect 52196 9432 52224 9608
rect 52730 9596 52736 9608
rect 52788 9596 52794 9648
rect 52914 9596 52920 9648
rect 52972 9636 52978 9648
rect 53101 9639 53159 9645
rect 53101 9636 53113 9639
rect 52972 9608 53113 9636
rect 52972 9596 52978 9608
rect 53101 9605 53113 9608
rect 53147 9605 53159 9639
rect 53101 9599 53159 9605
rect 53193 9639 53251 9645
rect 53193 9605 53205 9639
rect 53239 9636 53251 9639
rect 55769 9639 55827 9645
rect 53239 9608 53328 9636
rect 53239 9605 53251 9608
rect 53193 9599 53251 9605
rect 53300 9580 53328 9608
rect 55769 9605 55781 9639
rect 55815 9636 55827 9639
rect 56042 9636 56048 9648
rect 55815 9608 56048 9636
rect 55815 9605 55827 9608
rect 55769 9599 55827 9605
rect 52454 9528 52460 9580
rect 52512 9568 52518 9580
rect 53009 9571 53067 9577
rect 53009 9568 53021 9571
rect 52512 9540 53021 9568
rect 52512 9528 52518 9540
rect 53009 9537 53021 9540
rect 53055 9537 53067 9571
rect 53009 9531 53067 9537
rect 53282 9528 53288 9580
rect 53340 9528 53346 9580
rect 53377 9571 53435 9577
rect 53377 9537 53389 9571
rect 53423 9537 53435 9571
rect 53377 9531 53435 9537
rect 52365 9503 52423 9509
rect 52365 9469 52377 9503
rect 52411 9500 52423 9503
rect 52546 9500 52552 9512
rect 52411 9472 52552 9500
rect 52411 9469 52423 9472
rect 52365 9463 52423 9469
rect 52546 9460 52552 9472
rect 52604 9460 52610 9512
rect 52917 9503 52975 9509
rect 52917 9469 52929 9503
rect 52963 9469 52975 9503
rect 53392 9500 53420 9531
rect 53466 9528 53472 9580
rect 53524 9568 53530 9580
rect 53524 9540 53569 9568
rect 53524 9528 53530 9540
rect 53650 9528 53656 9580
rect 53708 9568 53714 9580
rect 54205 9571 54263 9577
rect 54205 9568 54217 9571
rect 53708 9540 54217 9568
rect 53708 9528 53714 9540
rect 54205 9537 54217 9540
rect 54251 9537 54263 9571
rect 54205 9531 54263 9537
rect 54447 9571 54505 9577
rect 54447 9537 54459 9571
rect 54493 9568 54505 9571
rect 55784 9568 55812 9599
rect 56042 9596 56048 9608
rect 56100 9596 56106 9648
rect 56428 9636 56456 9664
rect 56870 9636 56876 9648
rect 56428 9608 56876 9636
rect 56870 9596 56876 9608
rect 56928 9596 56934 9648
rect 58066 9636 58072 9648
rect 58027 9608 58072 9636
rect 58066 9596 58072 9608
rect 58124 9596 58130 9648
rect 56410 9568 56416 9580
rect 54493 9540 55812 9568
rect 56371 9540 56416 9568
rect 54493 9537 54505 9540
rect 54447 9531 54505 9537
rect 56410 9528 56416 9540
rect 56468 9528 56474 9580
rect 53742 9500 53748 9512
rect 53392 9472 53748 9500
rect 52917 9463 52975 9469
rect 49743 9404 52224 9432
rect 52273 9435 52331 9441
rect 49743 9401 49755 9404
rect 49697 9395 49755 9401
rect 52273 9401 52285 9435
rect 52319 9432 52331 9435
rect 52932 9432 52960 9463
rect 53742 9460 53748 9472
rect 53800 9460 53806 9512
rect 54570 9460 54576 9512
rect 54628 9500 54634 9512
rect 54757 9503 54815 9509
rect 54757 9500 54769 9503
rect 54628 9472 54769 9500
rect 54628 9460 54634 9472
rect 54757 9469 54769 9472
rect 54803 9469 54815 9503
rect 54757 9463 54815 9469
rect 54849 9503 54907 9509
rect 54849 9469 54861 9503
rect 54895 9500 54907 9503
rect 54895 9472 55536 9500
rect 54895 9469 54907 9472
rect 54849 9463 54907 9469
rect 55508 9444 55536 9472
rect 52319 9404 52960 9432
rect 52319 9401 52331 9404
rect 52273 9395 52331 9401
rect 47213 9367 47271 9373
rect 47213 9333 47225 9367
rect 47259 9364 47271 9367
rect 49712 9364 49740 9395
rect 53006 9392 53012 9444
rect 53064 9432 53070 9444
rect 55309 9435 55367 9441
rect 55309 9432 55321 9435
rect 53064 9404 55321 9432
rect 53064 9392 53070 9404
rect 55309 9401 55321 9404
rect 55355 9401 55367 9435
rect 55490 9432 55496 9444
rect 55451 9404 55496 9432
rect 55309 9395 55367 9401
rect 55490 9392 55496 9404
rect 55548 9392 55554 9444
rect 56870 9432 56876 9444
rect 56831 9404 56876 9432
rect 56870 9392 56876 9404
rect 56928 9392 56934 9444
rect 47259 9336 49740 9364
rect 47259 9333 47271 9336
rect 47213 9327 47271 9333
rect 49970 9324 49976 9376
rect 50028 9364 50034 9376
rect 50709 9367 50767 9373
rect 50709 9364 50721 9367
rect 50028 9336 50721 9364
rect 50028 9324 50034 9336
rect 50709 9333 50721 9336
rect 50755 9333 50767 9367
rect 50709 9327 50767 9333
rect 51074 9324 51080 9376
rect 51132 9364 51138 9376
rect 51353 9367 51411 9373
rect 51353 9364 51365 9367
rect 51132 9336 51365 9364
rect 51132 9324 51138 9336
rect 51353 9333 51365 9336
rect 51399 9364 51411 9367
rect 54018 9364 54024 9376
rect 51399 9336 54024 9364
rect 51399 9333 51411 9336
rect 51353 9327 51411 9333
rect 54018 9324 54024 9336
rect 54076 9364 54082 9376
rect 54846 9364 54852 9376
rect 54076 9336 54852 9364
rect 54076 9324 54082 9336
rect 54846 9324 54852 9336
rect 54904 9324 54910 9376
rect 56778 9324 56784 9376
rect 56836 9364 56842 9376
rect 57425 9367 57483 9373
rect 57425 9364 57437 9367
rect 56836 9336 57437 9364
rect 56836 9324 56842 9336
rect 57425 9333 57437 9336
rect 57471 9333 57483 9367
rect 57425 9327 57483 9333
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 26145 9163 26203 9169
rect 26145 9129 26157 9163
rect 26191 9160 26203 9163
rect 30377 9163 30435 9169
rect 30377 9160 30389 9163
rect 26191 9132 30389 9160
rect 26191 9129 26203 9132
rect 26145 9123 26203 9129
rect 30377 9129 30389 9132
rect 30423 9129 30435 9163
rect 30377 9123 30435 9129
rect 30745 9163 30803 9169
rect 30745 9129 30757 9163
rect 30791 9160 30803 9163
rect 30834 9160 30840 9172
rect 30791 9132 30840 9160
rect 30791 9129 30803 9132
rect 30745 9123 30803 9129
rect 25958 9052 25964 9104
rect 26016 9092 26022 9104
rect 26053 9095 26111 9101
rect 26053 9092 26065 9095
rect 26016 9064 26065 9092
rect 26016 9052 26022 9064
rect 26053 9061 26065 9064
rect 26099 9061 26111 9095
rect 26053 9055 26111 9061
rect 27525 9095 27583 9101
rect 27525 9061 27537 9095
rect 27571 9092 27583 9095
rect 27798 9092 27804 9104
rect 27571 9064 27804 9092
rect 27571 9061 27583 9064
rect 27525 9055 27583 9061
rect 27798 9052 27804 9064
rect 27856 9052 27862 9104
rect 28258 9092 28264 9104
rect 28000 9064 28264 9092
rect 24673 9027 24731 9033
rect 24673 8993 24685 9027
rect 24719 9024 24731 9027
rect 25225 9027 25283 9033
rect 25225 9024 25237 9027
rect 24719 8996 25237 9024
rect 24719 8993 24731 8996
rect 24673 8987 24731 8993
rect 25225 8993 25237 8996
rect 25271 9024 25283 9027
rect 25682 9024 25688 9036
rect 25271 8996 25688 9024
rect 25271 8993 25283 8996
rect 25225 8987 25283 8993
rect 25682 8984 25688 8996
rect 25740 9024 25746 9036
rect 28000 9033 28028 9064
rect 28258 9052 28264 9064
rect 28316 9052 28322 9104
rect 28902 9052 28908 9104
rect 28960 9092 28966 9104
rect 28997 9095 29055 9101
rect 28997 9092 29009 9095
rect 28960 9064 29009 9092
rect 28960 9052 28966 9064
rect 28997 9061 29009 9064
rect 29043 9061 29055 9095
rect 28997 9055 29055 9061
rect 29362 9052 29368 9104
rect 29420 9092 29426 9104
rect 29917 9095 29975 9101
rect 29917 9092 29929 9095
rect 29420 9064 29929 9092
rect 29420 9052 29426 9064
rect 29917 9061 29929 9064
rect 29963 9092 29975 9095
rect 30282 9092 30288 9104
rect 29963 9064 30288 9092
rect 29963 9061 29975 9064
rect 29917 9055 29975 9061
rect 30282 9052 30288 9064
rect 30340 9052 30346 9104
rect 30392 9092 30420 9123
rect 30834 9120 30840 9132
rect 30892 9120 30898 9172
rect 31570 9120 31576 9172
rect 31628 9160 31634 9172
rect 32401 9163 32459 9169
rect 32401 9160 32413 9163
rect 31628 9132 32413 9160
rect 31628 9120 31634 9132
rect 32401 9129 32413 9132
rect 32447 9129 32459 9163
rect 32401 9123 32459 9129
rect 32858 9120 32864 9172
rect 32916 9160 32922 9172
rect 32953 9163 33011 9169
rect 32953 9160 32965 9163
rect 32916 9132 32965 9160
rect 32916 9120 32922 9132
rect 32953 9129 32965 9132
rect 32999 9129 33011 9163
rect 32953 9123 33011 9129
rect 33042 9120 33048 9172
rect 33100 9160 33106 9172
rect 33413 9163 33471 9169
rect 33413 9160 33425 9163
rect 33100 9132 33425 9160
rect 33100 9120 33106 9132
rect 33413 9129 33425 9132
rect 33459 9129 33471 9163
rect 33413 9123 33471 9129
rect 33594 9120 33600 9172
rect 33652 9160 33658 9172
rect 33781 9163 33839 9169
rect 33781 9160 33793 9163
rect 33652 9132 33793 9160
rect 33652 9120 33658 9132
rect 33781 9129 33793 9132
rect 33827 9129 33839 9163
rect 33781 9123 33839 9129
rect 33870 9120 33876 9172
rect 33928 9160 33934 9172
rect 34790 9160 34796 9172
rect 33928 9132 34796 9160
rect 33928 9120 33934 9132
rect 34790 9120 34796 9132
rect 34848 9120 34854 9172
rect 35066 9120 35072 9172
rect 35124 9160 35130 9172
rect 35621 9163 35679 9169
rect 35621 9160 35633 9163
rect 35124 9132 35633 9160
rect 35124 9120 35130 9132
rect 35621 9129 35633 9132
rect 35667 9160 35679 9163
rect 35710 9160 35716 9172
rect 35667 9132 35716 9160
rect 35667 9129 35679 9132
rect 35621 9123 35679 9129
rect 35710 9120 35716 9132
rect 35768 9120 35774 9172
rect 36446 9120 36452 9172
rect 36504 9160 36510 9172
rect 37277 9163 37335 9169
rect 36504 9132 36860 9160
rect 36504 9120 36510 9132
rect 31481 9095 31539 9101
rect 31481 9092 31493 9095
rect 30392 9064 31493 9092
rect 31481 9061 31493 9064
rect 31527 9061 31539 9095
rect 31481 9055 31539 9061
rect 31754 9052 31760 9104
rect 31812 9092 31818 9104
rect 36722 9092 36728 9104
rect 31812 9064 36728 9092
rect 31812 9052 31818 9064
rect 36722 9052 36728 9064
rect 36780 9052 36786 9104
rect 36832 9092 36860 9132
rect 37277 9129 37289 9163
rect 37323 9160 37335 9163
rect 37458 9160 37464 9172
rect 37323 9132 37464 9160
rect 37323 9129 37335 9132
rect 37277 9123 37335 9129
rect 37458 9120 37464 9132
rect 37516 9120 37522 9172
rect 38378 9120 38384 9172
rect 38436 9160 38442 9172
rect 38657 9163 38715 9169
rect 38657 9160 38669 9163
rect 38436 9132 38669 9160
rect 38436 9120 38442 9132
rect 38657 9129 38669 9132
rect 38703 9129 38715 9163
rect 38838 9160 38844 9172
rect 38799 9132 38844 9160
rect 38657 9123 38715 9129
rect 38838 9120 38844 9132
rect 38896 9120 38902 9172
rect 39393 9163 39451 9169
rect 39393 9129 39405 9163
rect 39439 9160 39451 9163
rect 40678 9160 40684 9172
rect 39439 9132 40684 9160
rect 39439 9129 39451 9132
rect 39393 9123 39451 9129
rect 40678 9120 40684 9132
rect 40736 9120 40742 9172
rect 45649 9163 45707 9169
rect 45649 9129 45661 9163
rect 45695 9160 45707 9163
rect 46382 9160 46388 9172
rect 45695 9132 46388 9160
rect 45695 9129 45707 9132
rect 45649 9123 45707 9129
rect 46382 9120 46388 9132
rect 46440 9120 46446 9172
rect 49145 9163 49203 9169
rect 46492 9132 48314 9160
rect 37737 9095 37795 9101
rect 37737 9092 37749 9095
rect 36832 9064 37749 9092
rect 37737 9061 37749 9064
rect 37783 9061 37795 9095
rect 40586 9092 40592 9104
rect 37737 9055 37795 9061
rect 40236 9064 40592 9092
rect 27985 9027 28043 9033
rect 25740 8996 26464 9024
rect 25740 8984 25746 8996
rect 26068 8968 26096 8996
rect 25961 8959 26019 8965
rect 25961 8925 25973 8959
rect 26007 8925 26019 8959
rect 25961 8919 26019 8925
rect 25976 8888 26004 8919
rect 26050 8916 26056 8968
rect 26108 8916 26114 8968
rect 26436 8965 26464 8996
rect 27985 8993 27997 9027
rect 28031 8993 28043 9027
rect 29822 9024 29828 9036
rect 27985 8987 28043 8993
rect 28184 8996 29828 9024
rect 26237 8959 26295 8965
rect 26237 8925 26249 8959
rect 26283 8925 26295 8959
rect 26237 8919 26295 8925
rect 26421 8959 26479 8965
rect 26421 8925 26433 8959
rect 26467 8925 26479 8959
rect 26421 8919 26479 8925
rect 26252 8888 26280 8919
rect 26970 8916 26976 8968
rect 27028 8956 27034 8968
rect 27614 8956 27620 8968
rect 27028 8928 27620 8956
rect 27028 8916 27034 8928
rect 27614 8916 27620 8928
rect 27672 8956 27678 8968
rect 27709 8959 27767 8965
rect 27709 8956 27721 8959
rect 27672 8928 27721 8956
rect 27672 8916 27678 8928
rect 27709 8925 27721 8928
rect 27755 8925 27767 8959
rect 27890 8956 27896 8968
rect 27851 8928 27896 8956
rect 27709 8919 27767 8925
rect 27890 8916 27896 8928
rect 27948 8916 27954 8968
rect 28077 8959 28135 8965
rect 28077 8925 28089 8959
rect 28123 8956 28135 8959
rect 28184 8956 28212 8996
rect 29822 8984 29828 8996
rect 29880 8984 29886 9036
rect 30006 8984 30012 9036
rect 30064 9024 30070 9036
rect 30469 9027 30527 9033
rect 30469 9024 30481 9027
rect 30064 8996 30481 9024
rect 30064 8984 30070 8996
rect 30469 8993 30481 8996
rect 30515 9024 30527 9027
rect 31570 9024 31576 9036
rect 30515 8996 31576 9024
rect 30515 8993 30527 8996
rect 30469 8987 30527 8993
rect 31570 8984 31576 8996
rect 31628 8984 31634 9036
rect 32677 9027 32735 9033
rect 32677 8993 32689 9027
rect 32723 9024 32735 9027
rect 32723 8996 34652 9024
rect 32723 8993 32735 8996
rect 32677 8987 32735 8993
rect 34624 8968 34652 8996
rect 35250 8984 35256 9036
rect 35308 9024 35314 9036
rect 35308 8996 35848 9024
rect 35308 8984 35314 8996
rect 28123 8928 28212 8956
rect 28261 8959 28319 8965
rect 28123 8925 28135 8928
rect 28077 8919 28135 8925
rect 28261 8925 28273 8959
rect 28307 8956 28319 8959
rect 28994 8956 29000 8968
rect 28307 8928 29000 8956
rect 28307 8925 28319 8928
rect 28261 8919 28319 8925
rect 28994 8916 29000 8928
rect 29052 8916 29058 8968
rect 29086 8916 29092 8968
rect 29144 8956 29150 8968
rect 29181 8959 29239 8965
rect 29181 8956 29193 8959
rect 29144 8928 29193 8956
rect 29144 8916 29150 8928
rect 29181 8925 29193 8928
rect 29227 8925 29239 8959
rect 29181 8919 29239 8925
rect 29638 8916 29644 8968
rect 29696 8956 29702 8968
rect 29733 8959 29791 8965
rect 29733 8956 29745 8959
rect 29696 8928 29745 8956
rect 29696 8916 29702 8928
rect 29733 8925 29745 8928
rect 29779 8925 29791 8959
rect 29733 8919 29791 8925
rect 29917 8959 29975 8965
rect 29917 8925 29929 8959
rect 29963 8925 29975 8959
rect 30374 8956 30380 8968
rect 30335 8928 30380 8956
rect 29917 8919 29975 8925
rect 26510 8888 26516 8900
rect 25976 8860 26096 8888
rect 26252 8860 26516 8888
rect 24026 8820 24032 8832
rect 23987 8792 24032 8820
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 25590 8780 25596 8832
rect 25648 8820 25654 8832
rect 25685 8823 25743 8829
rect 25685 8820 25697 8823
rect 25648 8792 25697 8820
rect 25648 8780 25654 8792
rect 25685 8789 25697 8792
rect 25731 8789 25743 8823
rect 26068 8820 26096 8860
rect 26510 8848 26516 8860
rect 26568 8888 26574 8900
rect 26568 8860 27200 8888
rect 26568 8848 26574 8860
rect 26326 8820 26332 8832
rect 26068 8792 26332 8820
rect 25685 8783 25743 8789
rect 26326 8780 26332 8792
rect 26384 8780 26390 8832
rect 26786 8780 26792 8832
rect 26844 8820 26850 8832
rect 26973 8823 27031 8829
rect 26973 8820 26985 8823
rect 26844 8792 26985 8820
rect 26844 8780 26850 8792
rect 26973 8789 26985 8792
rect 27019 8789 27031 8823
rect 27172 8820 27200 8860
rect 27246 8848 27252 8900
rect 27304 8888 27310 8900
rect 28442 8888 28448 8900
rect 27304 8860 28448 8888
rect 27304 8848 27310 8860
rect 28442 8848 28448 8860
rect 28500 8888 28506 8900
rect 29546 8888 29552 8900
rect 28500 8860 29552 8888
rect 28500 8848 28506 8860
rect 29546 8848 29552 8860
rect 29604 8848 29610 8900
rect 29932 8888 29960 8919
rect 30374 8916 30380 8928
rect 30432 8956 30438 8968
rect 31386 8956 31392 8968
rect 30432 8928 31392 8956
rect 30432 8916 30438 8928
rect 31386 8916 31392 8928
rect 31444 8916 31450 8968
rect 31481 8959 31539 8965
rect 31481 8925 31493 8959
rect 31527 8925 31539 8959
rect 31481 8919 31539 8925
rect 31665 8959 31723 8965
rect 31665 8925 31677 8959
rect 31711 8956 31723 8959
rect 32769 8959 32827 8965
rect 31711 8928 32536 8956
rect 31711 8925 31723 8928
rect 31665 8919 31723 8925
rect 31496 8888 31524 8919
rect 32030 8888 32036 8900
rect 29932 8860 31432 8888
rect 31496 8860 32036 8888
rect 31404 8832 31432 8860
rect 32030 8848 32036 8860
rect 32088 8888 32094 8900
rect 32306 8888 32312 8900
rect 32088 8860 32168 8888
rect 32267 8860 32312 8888
rect 32088 8848 32094 8860
rect 30834 8820 30840 8832
rect 27172 8792 30840 8820
rect 26973 8783 27031 8789
rect 30834 8780 30840 8792
rect 30892 8780 30898 8832
rect 31386 8780 31392 8832
rect 31444 8780 31450 8832
rect 31662 8780 31668 8832
rect 31720 8820 31726 8832
rect 31846 8820 31852 8832
rect 31720 8792 31852 8820
rect 31720 8780 31726 8792
rect 31846 8780 31852 8792
rect 31904 8780 31910 8832
rect 32140 8820 32168 8860
rect 32306 8848 32312 8860
rect 32364 8848 32370 8900
rect 32214 8820 32220 8832
rect 32140 8792 32220 8820
rect 32214 8780 32220 8792
rect 32272 8780 32278 8832
rect 32508 8820 32536 8928
rect 32769 8925 32781 8959
rect 32815 8925 32827 8959
rect 32769 8919 32827 8925
rect 32784 8820 32812 8919
rect 32950 8916 32956 8968
rect 33008 8956 33014 8968
rect 33413 8959 33471 8965
rect 33413 8956 33425 8959
rect 33008 8928 33425 8956
rect 33008 8916 33014 8928
rect 33413 8925 33425 8928
rect 33459 8925 33471 8959
rect 33413 8919 33471 8925
rect 33594 8916 33600 8968
rect 33652 8956 33658 8968
rect 34146 8956 34152 8968
rect 33652 8928 34152 8956
rect 33652 8916 33658 8928
rect 34146 8916 34152 8928
rect 34204 8916 34210 8968
rect 34606 8916 34612 8968
rect 34664 8956 34670 8968
rect 34790 8956 34796 8968
rect 34664 8928 34796 8956
rect 34664 8916 34670 8928
rect 34790 8916 34796 8928
rect 34848 8956 34854 8968
rect 34885 8959 34943 8965
rect 34885 8956 34897 8959
rect 34848 8928 34897 8956
rect 34848 8916 34854 8928
rect 34885 8925 34897 8928
rect 34931 8925 34943 8959
rect 35066 8956 35072 8968
rect 35027 8928 35072 8956
rect 34885 8919 34943 8925
rect 35066 8916 35072 8928
rect 35124 8916 35130 8968
rect 35342 8916 35348 8968
rect 35400 8956 35406 8968
rect 35713 8959 35771 8965
rect 35713 8956 35725 8959
rect 35400 8928 35725 8956
rect 35400 8916 35406 8928
rect 35713 8925 35725 8928
rect 35759 8925 35771 8959
rect 35820 8956 35848 8996
rect 36630 8984 36636 9036
rect 36688 9024 36694 9036
rect 36817 9027 36875 9033
rect 36817 9024 36829 9027
rect 36688 8996 36829 9024
rect 36688 8984 36694 8996
rect 36817 8993 36829 8996
rect 36863 8993 36875 9027
rect 39574 9024 39580 9036
rect 36817 8987 36875 8993
rect 37016 8996 39580 9024
rect 36906 8956 36912 8968
rect 35820 8928 36912 8956
rect 35713 8919 35771 8925
rect 36906 8916 36912 8928
rect 36964 8916 36970 8968
rect 35084 8888 35112 8916
rect 33704 8860 35112 8888
rect 33704 8820 33732 8860
rect 35802 8848 35808 8900
rect 35860 8888 35866 8900
rect 36265 8891 36323 8897
rect 36265 8888 36277 8891
rect 35860 8860 36277 8888
rect 35860 8848 35866 8860
rect 36265 8857 36277 8860
rect 36311 8888 36323 8891
rect 37016 8888 37044 8996
rect 39574 8984 39580 8996
rect 39632 8984 39638 9036
rect 37090 8916 37096 8968
rect 37148 8956 37154 8968
rect 38473 8959 38531 8965
rect 38473 8956 38485 8959
rect 37148 8928 38485 8956
rect 37148 8916 37154 8928
rect 38473 8925 38485 8928
rect 38519 8925 38531 8959
rect 38473 8919 38531 8925
rect 38749 8959 38807 8965
rect 38749 8925 38761 8959
rect 38795 8956 38807 8959
rect 38930 8956 38936 8968
rect 38795 8928 38936 8956
rect 38795 8925 38807 8928
rect 38749 8919 38807 8925
rect 38930 8916 38936 8928
rect 38988 8916 38994 8968
rect 40236 8965 40264 9064
rect 40586 9052 40592 9064
rect 40644 9092 40650 9104
rect 41233 9095 41291 9101
rect 41233 9092 41245 9095
rect 40644 9064 41245 9092
rect 40644 9052 40650 9064
rect 41233 9061 41245 9064
rect 41279 9061 41291 9095
rect 41233 9055 41291 9061
rect 42429 9095 42487 9101
rect 42429 9061 42441 9095
rect 42475 9092 42487 9095
rect 42518 9092 42524 9104
rect 42475 9064 42524 9092
rect 42475 9061 42487 9064
rect 42429 9055 42487 9061
rect 42518 9052 42524 9064
rect 42576 9052 42582 9104
rect 42794 9052 42800 9104
rect 42852 9092 42858 9104
rect 43530 9092 43536 9104
rect 42852 9064 43536 9092
rect 42852 9052 42858 9064
rect 43530 9052 43536 9064
rect 43588 9092 43594 9104
rect 45094 9092 45100 9104
rect 43588 9064 45100 9092
rect 43588 9052 43594 9064
rect 45094 9052 45100 9064
rect 45152 9092 45158 9104
rect 46492 9092 46520 9132
rect 45152 9064 46520 9092
rect 45152 9052 45158 9064
rect 47026 9052 47032 9104
rect 47084 9092 47090 9104
rect 48286 9092 48314 9132
rect 49145 9129 49157 9163
rect 49191 9160 49203 9163
rect 50246 9160 50252 9172
rect 49191 9132 50252 9160
rect 49191 9129 49203 9132
rect 49145 9123 49203 9129
rect 50246 9120 50252 9132
rect 50304 9120 50310 9172
rect 50798 9160 50804 9172
rect 50759 9132 50804 9160
rect 50798 9120 50804 9132
rect 50856 9120 50862 9172
rect 53193 9163 53251 9169
rect 53193 9129 53205 9163
rect 53239 9160 53251 9163
rect 54202 9160 54208 9172
rect 53239 9132 54208 9160
rect 53239 9129 53251 9132
rect 53193 9123 53251 9129
rect 54202 9120 54208 9132
rect 54260 9120 54266 9172
rect 55585 9163 55643 9169
rect 55585 9129 55597 9163
rect 55631 9160 55643 9163
rect 55674 9160 55680 9172
rect 55631 9132 55680 9160
rect 55631 9129 55643 9132
rect 55585 9123 55643 9129
rect 55674 9120 55680 9132
rect 55732 9120 55738 9172
rect 56137 9163 56195 9169
rect 56137 9129 56149 9163
rect 56183 9160 56195 9163
rect 56594 9160 56600 9172
rect 56183 9132 56600 9160
rect 56183 9129 56195 9132
rect 56137 9123 56195 9129
rect 56594 9120 56600 9132
rect 56652 9120 56658 9172
rect 49602 9092 49608 9104
rect 47084 9064 47129 9092
rect 48286 9064 49608 9092
rect 47084 9052 47090 9064
rect 49602 9052 49608 9064
rect 49660 9052 49666 9104
rect 49786 9052 49792 9104
rect 49844 9092 49850 9104
rect 50893 9095 50951 9101
rect 50893 9092 50905 9095
rect 49844 9064 50905 9092
rect 49844 9052 49850 9064
rect 50893 9061 50905 9064
rect 50939 9092 50951 9095
rect 51350 9092 51356 9104
rect 50939 9064 51356 9092
rect 50939 9061 50951 9064
rect 50893 9055 50951 9061
rect 51350 9052 51356 9064
rect 51408 9052 51414 9104
rect 51534 9052 51540 9104
rect 51592 9092 51598 9104
rect 51721 9095 51779 9101
rect 51721 9092 51733 9095
rect 51592 9064 51733 9092
rect 51592 9052 51598 9064
rect 51721 9061 51733 9064
rect 51767 9061 51779 9095
rect 51721 9055 51779 9061
rect 51828 9064 54248 9092
rect 40402 8984 40408 9036
rect 40460 9024 40466 9036
rect 41322 9024 41328 9036
rect 40460 8996 40632 9024
rect 41283 8996 41328 9024
rect 40460 8984 40466 8996
rect 40604 8965 40632 8996
rect 41322 8984 41328 8996
rect 41380 8984 41386 9036
rect 42812 9024 42840 9052
rect 42076 8996 42840 9024
rect 40221 8959 40279 8965
rect 40221 8925 40233 8959
rect 40267 8925 40279 8959
rect 40221 8919 40279 8925
rect 40589 8959 40647 8965
rect 40589 8925 40601 8959
rect 40635 8925 40647 8959
rect 41046 8956 41052 8968
rect 41007 8928 41052 8956
rect 40589 8919 40647 8925
rect 41046 8916 41052 8928
rect 41104 8916 41110 8968
rect 41138 8916 41144 8968
rect 41196 8956 41202 8968
rect 41196 8928 41241 8956
rect 41196 8916 41202 8928
rect 41782 8916 41788 8968
rect 41840 8956 41846 8968
rect 42076 8965 42104 8996
rect 43622 8984 43628 9036
rect 43680 9024 43686 9036
rect 44910 9024 44916 9036
rect 43680 8996 44916 9024
rect 43680 8984 43686 8996
rect 44910 8984 44916 8996
rect 44968 8984 44974 9036
rect 45922 8984 45928 9036
rect 45980 8984 45986 9036
rect 46014 8984 46020 9036
rect 46072 9024 46078 9036
rect 46072 8996 46796 9024
rect 46072 8984 46078 8996
rect 42061 8959 42119 8965
rect 42061 8956 42073 8959
rect 41840 8928 42073 8956
rect 41840 8916 41846 8928
rect 42061 8925 42073 8928
rect 42107 8925 42119 8959
rect 42061 8919 42119 8925
rect 42150 8916 42156 8968
rect 42208 8956 42214 8968
rect 44818 8956 44824 8968
rect 42208 8928 42253 8956
rect 44192 8928 44824 8956
rect 42208 8916 42214 8928
rect 38378 8888 38384 8900
rect 36311 8860 37044 8888
rect 38339 8860 38384 8888
rect 36311 8857 36323 8860
rect 36265 8851 36323 8857
rect 38378 8848 38384 8860
rect 38436 8848 38442 8900
rect 39758 8848 39764 8900
rect 39816 8888 39822 8900
rect 40313 8891 40371 8897
rect 40313 8888 40325 8891
rect 39816 8860 40325 8888
rect 39816 8848 39822 8860
rect 40313 8857 40325 8860
rect 40359 8857 40371 8891
rect 40313 8851 40371 8857
rect 40402 8848 40408 8900
rect 40460 8888 40466 8900
rect 42981 8891 43039 8897
rect 40460 8860 40505 8888
rect 40460 8848 40466 8860
rect 42981 8857 42993 8891
rect 43027 8888 43039 8891
rect 43438 8888 43444 8900
rect 43027 8860 43444 8888
rect 43027 8857 43039 8860
rect 42981 8851 43039 8857
rect 43438 8848 43444 8860
rect 43496 8848 43502 8900
rect 43622 8848 43628 8900
rect 43680 8888 43686 8900
rect 44192 8897 44220 8928
rect 44818 8916 44824 8928
rect 44876 8916 44882 8968
rect 45278 8916 45284 8968
rect 45336 8956 45342 8968
rect 45833 8959 45891 8965
rect 45336 8928 45787 8956
rect 45336 8916 45342 8928
rect 44177 8891 44235 8897
rect 44177 8888 44189 8891
rect 43680 8860 44189 8888
rect 43680 8848 43686 8860
rect 44177 8857 44189 8860
rect 44223 8857 44235 8891
rect 44177 8851 44235 8857
rect 44545 8891 44603 8897
rect 44545 8857 44557 8891
rect 44591 8888 44603 8891
rect 45554 8888 45560 8900
rect 44591 8860 45560 8888
rect 44591 8857 44603 8860
rect 44545 8851 44603 8857
rect 45554 8848 45560 8860
rect 45612 8848 45618 8900
rect 45759 8888 45787 8928
rect 45833 8925 45845 8959
rect 45879 8956 45891 8959
rect 45940 8956 45968 8984
rect 46106 8956 46112 8968
rect 45879 8928 45968 8956
rect 46067 8928 46112 8956
rect 45879 8925 45891 8928
rect 45833 8919 45891 8925
rect 46106 8916 46112 8928
rect 46164 8916 46170 8968
rect 46290 8956 46296 8968
rect 46251 8928 46296 8956
rect 46290 8916 46296 8928
rect 46348 8916 46354 8968
rect 46768 8965 46796 8996
rect 46952 8996 48636 9024
rect 46753 8959 46811 8965
rect 46753 8925 46765 8959
rect 46799 8925 46811 8959
rect 46753 8919 46811 8925
rect 45925 8891 45983 8897
rect 45925 8888 45937 8891
rect 45759 8860 45937 8888
rect 45925 8857 45937 8860
rect 45971 8857 45983 8891
rect 45925 8851 45983 8857
rect 46017 8891 46075 8897
rect 46017 8857 46029 8891
rect 46063 8857 46075 8891
rect 46017 8851 46075 8857
rect 34330 8820 34336 8832
rect 32508 8792 33732 8820
rect 34291 8792 34336 8820
rect 34330 8780 34336 8792
rect 34388 8780 34394 8832
rect 34974 8820 34980 8832
rect 34935 8792 34980 8820
rect 34974 8780 34980 8792
rect 35032 8780 35038 8832
rect 35986 8780 35992 8832
rect 36044 8820 36050 8832
rect 37458 8820 37464 8832
rect 36044 8792 37464 8820
rect 36044 8780 36050 8792
rect 37458 8780 37464 8792
rect 37516 8780 37522 8832
rect 40037 8823 40095 8829
rect 40037 8789 40049 8823
rect 40083 8820 40095 8823
rect 40126 8820 40132 8832
rect 40083 8792 40132 8820
rect 40083 8789 40095 8792
rect 40037 8783 40095 8789
rect 40126 8780 40132 8792
rect 40184 8780 40190 8832
rect 43162 8780 43168 8832
rect 43220 8820 43226 8832
rect 43533 8823 43591 8829
rect 43533 8820 43545 8823
rect 43220 8792 43545 8820
rect 43220 8780 43226 8792
rect 43533 8789 43545 8792
rect 43579 8820 43591 8823
rect 44082 8820 44088 8832
rect 43579 8792 44088 8820
rect 43579 8789 43591 8792
rect 43533 8783 43591 8789
rect 44082 8780 44088 8792
rect 44140 8820 44146 8832
rect 44634 8820 44640 8832
rect 44140 8792 44640 8820
rect 44140 8780 44146 8792
rect 44634 8780 44640 8792
rect 44692 8780 44698 8832
rect 46032 8820 46060 8851
rect 46198 8848 46204 8900
rect 46256 8888 46262 8900
rect 46845 8891 46903 8897
rect 46845 8888 46857 8891
rect 46256 8860 46857 8888
rect 46256 8848 46262 8860
rect 46845 8857 46857 8860
rect 46891 8857 46903 8891
rect 46845 8851 46903 8857
rect 46566 8820 46572 8832
rect 46032 8792 46572 8820
rect 46566 8780 46572 8792
rect 46624 8820 46630 8832
rect 46952 8820 46980 8996
rect 47210 8916 47216 8968
rect 47268 8956 47274 8968
rect 47673 8959 47731 8965
rect 47673 8956 47685 8959
rect 47268 8928 47685 8956
rect 47268 8916 47274 8928
rect 47673 8925 47685 8928
rect 47719 8925 47731 8959
rect 48498 8956 48504 8968
rect 47673 8919 47731 8925
rect 48148 8928 48504 8956
rect 47029 8891 47087 8897
rect 47029 8857 47041 8891
rect 47075 8888 47087 8891
rect 48148 8888 48176 8928
rect 48498 8916 48504 8928
rect 48556 8916 48562 8968
rect 48608 8965 48636 8996
rect 50062 8984 50068 9036
rect 50120 9024 50126 9036
rect 51828 9024 51856 9064
rect 52546 9024 52552 9036
rect 50120 8996 51856 9024
rect 51920 8996 52552 9024
rect 50120 8984 50126 8996
rect 48593 8959 48651 8965
rect 48593 8925 48605 8959
rect 48639 8956 48651 8959
rect 49234 8956 49240 8968
rect 48639 8928 49240 8956
rect 48639 8925 48651 8928
rect 48593 8919 48651 8925
rect 49234 8916 49240 8928
rect 49292 8916 49298 8968
rect 49970 8916 49976 8968
rect 50028 8956 50034 8968
rect 51920 8965 51948 8996
rect 52546 8984 52552 8996
rect 52604 8984 52610 9036
rect 53926 9024 53932 9036
rect 53887 8996 53932 9024
rect 53926 8984 53932 8996
rect 53984 8984 53990 9036
rect 54018 8984 54024 9036
rect 54076 9024 54082 9036
rect 54220 9024 54248 9064
rect 54478 9052 54484 9104
rect 54536 9092 54542 9104
rect 54849 9095 54907 9101
rect 54849 9092 54861 9095
rect 54536 9064 54861 9092
rect 54536 9052 54542 9064
rect 54849 9061 54861 9064
rect 54895 9092 54907 9095
rect 56318 9092 56324 9104
rect 54895 9064 56324 9092
rect 54895 9061 54907 9064
rect 54849 9055 54907 9061
rect 56318 9052 56324 9064
rect 56376 9052 56382 9104
rect 58253 9095 58311 9101
rect 58253 9092 58265 9095
rect 57946 9064 58265 9092
rect 55398 9024 55404 9036
rect 54076 8996 54121 9024
rect 54220 8996 55404 9024
rect 54076 8984 54082 8996
rect 51905 8959 51963 8965
rect 50028 8928 51856 8956
rect 50028 8916 50034 8928
rect 47075 8860 48176 8888
rect 48225 8891 48283 8897
rect 47075 8857 47087 8860
rect 47029 8851 47087 8857
rect 48225 8857 48237 8891
rect 48271 8857 48283 8891
rect 48225 8851 48283 8857
rect 47578 8820 47584 8832
rect 46624 8792 46980 8820
rect 47539 8792 47584 8820
rect 46624 8780 46630 8792
rect 47578 8780 47584 8792
rect 47636 8780 47642 8832
rect 47762 8780 47768 8832
rect 47820 8820 47826 8832
rect 48130 8820 48136 8832
rect 47820 8792 48136 8820
rect 47820 8780 47826 8792
rect 48130 8780 48136 8792
rect 48188 8820 48194 8832
rect 48240 8820 48268 8851
rect 49602 8848 49608 8900
rect 49660 8888 49666 8900
rect 51261 8891 51319 8897
rect 51261 8888 51273 8891
rect 49660 8860 51273 8888
rect 49660 8848 49666 8860
rect 51261 8857 51273 8860
rect 51307 8888 51319 8891
rect 51718 8888 51724 8900
rect 51307 8860 51724 8888
rect 51307 8857 51319 8860
rect 51261 8851 51319 8857
rect 51718 8848 51724 8860
rect 51776 8848 51782 8900
rect 51828 8888 51856 8928
rect 51905 8925 51917 8959
rect 51951 8925 51963 8959
rect 51905 8919 51963 8925
rect 52012 8928 52592 8956
rect 52012 8888 52040 8928
rect 51828 8860 52040 8888
rect 52089 8891 52147 8897
rect 52089 8857 52101 8891
rect 52135 8857 52147 8891
rect 52564 8888 52592 8928
rect 52638 8916 52644 8968
rect 52696 8956 52702 8968
rect 53009 8959 53067 8965
rect 53009 8956 53021 8959
rect 52696 8928 53021 8956
rect 52696 8916 52702 8928
rect 53009 8925 53021 8928
rect 53055 8925 53067 8959
rect 53009 8919 53067 8925
rect 53193 8959 53251 8965
rect 53193 8925 53205 8959
rect 53239 8956 53251 8959
rect 53653 8959 53711 8965
rect 53653 8956 53665 8959
rect 53239 8928 53665 8956
rect 53239 8925 53251 8928
rect 53193 8919 53251 8925
rect 53653 8925 53665 8928
rect 53699 8925 53711 8959
rect 53653 8919 53711 8925
rect 53837 8959 53895 8965
rect 53837 8925 53849 8959
rect 53883 8925 53895 8959
rect 53837 8919 53895 8925
rect 54113 8959 54171 8965
rect 54113 8925 54125 8959
rect 54159 8956 54171 8959
rect 54220 8956 54248 8996
rect 55398 8984 55404 8996
rect 55456 8984 55462 9036
rect 54159 8928 54248 8956
rect 54297 8959 54355 8965
rect 54159 8925 54171 8928
rect 54113 8919 54171 8925
rect 54297 8925 54309 8959
rect 54343 8956 54355 8959
rect 54386 8956 54392 8968
rect 54343 8928 54392 8956
rect 54343 8925 54355 8928
rect 54297 8919 54355 8925
rect 52730 8888 52736 8900
rect 52564 8860 52736 8888
rect 52089 8851 52147 8857
rect 48188 8792 48268 8820
rect 48188 8780 48194 8792
rect 48314 8780 48320 8832
rect 48372 8820 48378 8832
rect 49142 8820 49148 8832
rect 48372 8792 49148 8820
rect 48372 8780 48378 8792
rect 49142 8780 49148 8792
rect 49200 8820 49206 8832
rect 49697 8823 49755 8829
rect 49697 8820 49709 8823
rect 49200 8792 49709 8820
rect 49200 8780 49206 8792
rect 49697 8789 49709 8792
rect 49743 8820 49755 8823
rect 50890 8820 50896 8832
rect 49743 8792 50896 8820
rect 49743 8789 49755 8792
rect 49697 8783 49755 8789
rect 50890 8780 50896 8792
rect 50948 8780 50954 8832
rect 51166 8780 51172 8832
rect 51224 8820 51230 8832
rect 52104 8820 52132 8851
rect 52730 8848 52736 8860
rect 52788 8888 52794 8900
rect 53852 8888 53880 8919
rect 54386 8916 54392 8928
rect 54444 8916 54450 8968
rect 56502 8916 56508 8968
rect 56560 8956 56566 8968
rect 57149 8959 57207 8965
rect 57149 8956 57161 8959
rect 56560 8928 57161 8956
rect 56560 8916 56566 8928
rect 57149 8925 57161 8928
rect 57195 8956 57207 8959
rect 57946 8956 57974 9064
rect 58253 9061 58265 9064
rect 58299 9061 58311 9095
rect 58253 9055 58311 9061
rect 57195 8928 57974 8956
rect 57195 8925 57207 8928
rect 57149 8919 57207 8925
rect 57330 8888 57336 8900
rect 52788 8860 57336 8888
rect 52788 8848 52794 8860
rect 57330 8848 57336 8860
rect 57388 8848 57394 8900
rect 51224 8792 52132 8820
rect 51224 8780 51230 8792
rect 53006 8780 53012 8832
rect 53064 8820 53070 8832
rect 54570 8820 54576 8832
rect 53064 8792 54576 8820
rect 53064 8780 53070 8792
rect 54570 8780 54576 8792
rect 54628 8780 54634 8832
rect 56686 8820 56692 8832
rect 56647 8792 56692 8820
rect 56686 8780 56692 8792
rect 56744 8780 56750 8832
rect 56870 8780 56876 8832
rect 56928 8820 56934 8832
rect 57701 8823 57759 8829
rect 57701 8820 57713 8823
rect 56928 8792 57713 8820
rect 56928 8780 56934 8792
rect 57701 8789 57713 8792
rect 57747 8789 57759 8823
rect 57701 8783 57759 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 25041 8619 25099 8625
rect 25041 8585 25053 8619
rect 25087 8616 25099 8619
rect 25314 8616 25320 8628
rect 25087 8588 25320 8616
rect 25087 8585 25099 8588
rect 25041 8579 25099 8585
rect 25314 8576 25320 8588
rect 25372 8576 25378 8628
rect 26694 8576 26700 8628
rect 26752 8616 26758 8628
rect 27801 8619 27859 8625
rect 27801 8616 27813 8619
rect 26752 8588 27813 8616
rect 26752 8576 26758 8588
rect 27801 8585 27813 8588
rect 27847 8585 27859 8619
rect 27801 8579 27859 8585
rect 28626 8576 28632 8628
rect 28684 8616 28690 8628
rect 28721 8619 28779 8625
rect 28721 8616 28733 8619
rect 28684 8588 28733 8616
rect 28684 8576 28690 8588
rect 28721 8585 28733 8588
rect 28767 8585 28779 8619
rect 28721 8579 28779 8585
rect 28828 8588 30420 8616
rect 25590 8548 25596 8560
rect 25551 8520 25596 8548
rect 25590 8508 25596 8520
rect 25648 8508 25654 8560
rect 25685 8551 25743 8557
rect 25685 8517 25697 8551
rect 25731 8548 25743 8551
rect 25866 8548 25872 8560
rect 25731 8520 25872 8548
rect 25731 8517 25743 8520
rect 25685 8511 25743 8517
rect 25866 8508 25872 8520
rect 25924 8508 25930 8560
rect 26602 8548 26608 8560
rect 26515 8520 26608 8548
rect 26602 8508 26608 8520
rect 26660 8548 26666 8560
rect 26660 8520 27568 8548
rect 26660 8508 26666 8520
rect 25314 8480 25320 8492
rect 25275 8452 25320 8480
rect 25314 8440 25320 8452
rect 25372 8440 25378 8492
rect 27154 8480 27160 8492
rect 27115 8452 27160 8480
rect 27154 8440 27160 8452
rect 27212 8440 27218 8492
rect 27540 8480 27568 8520
rect 28258 8508 28264 8560
rect 28316 8548 28322 8560
rect 28828 8548 28856 8588
rect 28316 8520 28856 8548
rect 29825 8551 29883 8557
rect 28316 8508 28322 8520
rect 29825 8517 29837 8551
rect 29871 8548 29883 8551
rect 30190 8548 30196 8560
rect 29871 8520 30196 8548
rect 29871 8517 29883 8520
rect 29825 8511 29883 8517
rect 30190 8508 30196 8520
rect 30248 8508 30254 8560
rect 27613 8483 27671 8489
rect 27613 8480 27625 8483
rect 27540 8452 27625 8480
rect 27613 8449 27625 8452
rect 27659 8449 27671 8483
rect 27613 8443 27671 8449
rect 28442 8440 28448 8492
rect 28500 8480 28506 8492
rect 28626 8480 28632 8492
rect 28500 8452 28632 8480
rect 28500 8440 28506 8452
rect 28626 8440 28632 8452
rect 28684 8480 28690 8492
rect 28905 8483 28963 8489
rect 28905 8480 28917 8483
rect 28684 8452 28917 8480
rect 28684 8440 28690 8452
rect 28905 8449 28917 8452
rect 28951 8449 28963 8483
rect 28905 8443 28963 8449
rect 29181 8483 29239 8489
rect 29181 8449 29193 8483
rect 29227 8480 29239 8483
rect 29270 8480 29276 8492
rect 29227 8452 29276 8480
rect 29227 8449 29239 8452
rect 29181 8443 29239 8449
rect 29270 8440 29276 8452
rect 29328 8440 29334 8492
rect 29546 8440 29552 8492
rect 29604 8480 29610 8492
rect 29733 8483 29791 8489
rect 29733 8480 29745 8483
rect 29604 8452 29745 8480
rect 29604 8440 29610 8452
rect 29733 8449 29745 8452
rect 29779 8449 29791 8483
rect 29733 8443 29791 8449
rect 29917 8483 29975 8489
rect 29917 8449 29929 8483
rect 29963 8480 29975 8483
rect 30006 8480 30012 8492
rect 29963 8452 30012 8480
rect 29963 8449 29975 8452
rect 29917 8443 29975 8449
rect 30006 8440 30012 8452
rect 30064 8440 30070 8492
rect 30392 8480 30420 8588
rect 31294 8576 31300 8628
rect 31352 8616 31358 8628
rect 32677 8619 32735 8625
rect 32677 8616 32689 8619
rect 31352 8588 32689 8616
rect 31352 8576 31358 8588
rect 32677 8585 32689 8588
rect 32723 8616 32735 8619
rect 37090 8616 37096 8628
rect 32723 8588 37096 8616
rect 32723 8585 32735 8588
rect 32677 8579 32735 8585
rect 37090 8576 37096 8588
rect 37148 8576 37154 8628
rect 37550 8616 37556 8628
rect 37511 8588 37556 8616
rect 37550 8576 37556 8588
rect 37608 8576 37614 8628
rect 38930 8616 38936 8628
rect 38891 8588 38936 8616
rect 38930 8576 38936 8588
rect 38988 8576 38994 8628
rect 43990 8616 43996 8628
rect 43951 8588 43996 8616
rect 43990 8576 43996 8588
rect 44048 8576 44054 8628
rect 46106 8576 46112 8628
rect 46164 8616 46170 8628
rect 47857 8619 47915 8625
rect 47857 8616 47869 8619
rect 46164 8588 47869 8616
rect 46164 8576 46170 8588
rect 47857 8585 47869 8588
rect 47903 8585 47915 8619
rect 47857 8579 47915 8585
rect 48314 8576 48320 8628
rect 48372 8616 48378 8628
rect 48777 8619 48835 8625
rect 48777 8616 48789 8619
rect 48372 8588 48789 8616
rect 48372 8576 48378 8588
rect 48777 8585 48789 8588
rect 48823 8616 48835 8619
rect 49786 8616 49792 8628
rect 48823 8588 49792 8616
rect 48823 8585 48835 8588
rect 48777 8579 48835 8585
rect 49786 8576 49792 8588
rect 49844 8576 49850 8628
rect 50706 8616 50712 8628
rect 50667 8588 50712 8616
rect 50706 8576 50712 8588
rect 50764 8576 50770 8628
rect 51350 8576 51356 8628
rect 51408 8616 51414 8628
rect 53006 8616 53012 8628
rect 51408 8588 53012 8616
rect 51408 8576 51414 8588
rect 53006 8576 53012 8588
rect 53064 8576 53070 8628
rect 53190 8576 53196 8628
rect 53248 8616 53254 8628
rect 54018 8616 54024 8628
rect 53248 8588 54024 8616
rect 53248 8576 53254 8588
rect 54018 8576 54024 8588
rect 54076 8576 54082 8628
rect 54662 8616 54668 8628
rect 54623 8588 54668 8616
rect 54662 8576 54668 8588
rect 54720 8576 54726 8628
rect 54846 8576 54852 8628
rect 54904 8616 54910 8628
rect 55306 8616 55312 8628
rect 54904 8588 55312 8616
rect 54904 8576 54910 8588
rect 55306 8576 55312 8588
rect 55364 8576 55370 8628
rect 56686 8576 56692 8628
rect 56744 8616 56750 8628
rect 58069 8619 58127 8625
rect 58069 8616 58081 8619
rect 56744 8588 58081 8616
rect 56744 8576 56750 8588
rect 58069 8585 58081 8588
rect 58115 8585 58127 8619
rect 58069 8579 58127 8585
rect 30466 8508 30472 8560
rect 30524 8548 30530 8560
rect 30745 8551 30803 8557
rect 30745 8548 30757 8551
rect 30524 8520 30757 8548
rect 30524 8508 30530 8520
rect 30745 8517 30757 8520
rect 30791 8517 30803 8551
rect 32490 8548 32496 8560
rect 30745 8511 30803 8517
rect 30944 8520 32496 8548
rect 30944 8489 30972 8520
rect 32490 8508 32496 8520
rect 32548 8548 32554 8560
rect 32858 8548 32864 8560
rect 32548 8520 32864 8548
rect 32548 8508 32554 8520
rect 32858 8508 32864 8520
rect 32916 8508 32922 8560
rect 34974 8548 34980 8560
rect 33888 8520 34980 8548
rect 30561 8483 30619 8489
rect 30561 8480 30573 8483
rect 30392 8452 30573 8480
rect 30561 8449 30573 8452
rect 30607 8449 30619 8483
rect 30561 8443 30619 8449
rect 30929 8483 30987 8489
rect 30929 8449 30941 8483
rect 30975 8449 30987 8483
rect 30929 8443 30987 8449
rect 31205 8483 31263 8489
rect 31205 8449 31217 8483
rect 31251 8480 31263 8483
rect 31386 8480 31392 8492
rect 31251 8452 31392 8480
rect 31251 8449 31263 8452
rect 31205 8443 31263 8449
rect 31386 8440 31392 8452
rect 31444 8440 31450 8492
rect 31757 8483 31815 8489
rect 31757 8449 31769 8483
rect 31803 8480 31815 8483
rect 31846 8480 31852 8492
rect 31803 8452 31852 8480
rect 31803 8449 31815 8452
rect 31757 8443 31815 8449
rect 31846 8440 31852 8452
rect 31904 8440 31910 8492
rect 32677 8483 32735 8489
rect 32677 8449 32689 8483
rect 32723 8480 32735 8483
rect 33226 8480 33232 8492
rect 32723 8452 33232 8480
rect 32723 8449 32735 8452
rect 32677 8443 32735 8449
rect 33226 8440 33232 8452
rect 33284 8480 33290 8492
rect 33594 8480 33600 8492
rect 33284 8452 33600 8480
rect 33284 8440 33290 8452
rect 33594 8440 33600 8452
rect 33652 8440 33658 8492
rect 33888 8489 33916 8520
rect 34974 8508 34980 8520
rect 35032 8508 35038 8560
rect 35710 8508 35716 8560
rect 35768 8548 35774 8560
rect 37568 8548 37596 8576
rect 35768 8520 36492 8548
rect 35768 8508 35774 8520
rect 33853 8483 33916 8489
rect 33853 8449 33865 8483
rect 33899 8450 33916 8483
rect 33965 8483 34023 8489
rect 33899 8449 33911 8450
rect 33853 8443 33911 8449
rect 33965 8449 33977 8483
rect 34011 8449 34023 8483
rect 33965 8443 34023 8449
rect 34062 8483 34120 8489
rect 34062 8449 34074 8483
rect 34108 8480 34120 8483
rect 34241 8483 34299 8489
rect 34108 8452 34192 8480
rect 34108 8449 34120 8452
rect 34062 8443 34120 8449
rect 23937 8415 23995 8421
rect 23937 8381 23949 8415
rect 23983 8412 23995 8415
rect 24026 8412 24032 8424
rect 23983 8384 24032 8412
rect 23983 8381 23995 8384
rect 23937 8375 23995 8381
rect 24026 8372 24032 8384
rect 24084 8412 24090 8424
rect 24489 8415 24547 8421
rect 24489 8412 24501 8415
rect 24084 8384 24501 8412
rect 24084 8372 24090 8384
rect 24489 8381 24501 8384
rect 24535 8412 24547 8415
rect 25205 8415 25263 8421
rect 25205 8412 25217 8415
rect 24535 8384 25217 8412
rect 24535 8381 24547 8384
rect 24489 8375 24547 8381
rect 25205 8381 25217 8384
rect 25251 8412 25263 8415
rect 26326 8412 26332 8424
rect 25251 8384 26332 8412
rect 25251 8381 25263 8384
rect 25205 8375 25263 8381
rect 26326 8372 26332 8384
rect 26384 8412 26390 8424
rect 27341 8415 27399 8421
rect 27341 8412 27353 8415
rect 26384 8384 27353 8412
rect 26384 8372 26390 8384
rect 27341 8381 27353 8384
rect 27387 8381 27399 8415
rect 27341 8375 27399 8381
rect 27430 8372 27436 8424
rect 27488 8412 27494 8424
rect 28997 8415 29055 8421
rect 27488 8384 27533 8412
rect 27488 8372 27494 8384
rect 28997 8381 29009 8415
rect 29043 8412 29055 8415
rect 30282 8412 30288 8424
rect 29043 8384 30288 8412
rect 29043 8381 29055 8384
rect 28997 8375 29055 8381
rect 30282 8372 30288 8384
rect 30340 8372 30346 8424
rect 30377 8415 30435 8421
rect 30377 8381 30389 8415
rect 30423 8412 30435 8415
rect 30466 8412 30472 8424
rect 30423 8384 30472 8412
rect 30423 8381 30435 8384
rect 30377 8375 30435 8381
rect 30466 8372 30472 8384
rect 30524 8372 30530 8424
rect 30834 8372 30840 8424
rect 30892 8412 30898 8424
rect 32309 8415 32367 8421
rect 32309 8412 32321 8415
rect 30892 8384 32321 8412
rect 30892 8372 30898 8384
rect 32309 8381 32321 8384
rect 32355 8412 32367 8415
rect 32766 8412 32772 8424
rect 32355 8384 32772 8412
rect 32355 8381 32367 8384
rect 32309 8375 32367 8381
rect 32766 8372 32772 8384
rect 32824 8372 32830 8424
rect 32858 8372 32864 8424
rect 32916 8412 32922 8424
rect 32916 8384 32961 8412
rect 32916 8372 32922 8384
rect 33686 8372 33692 8424
rect 33744 8412 33750 8424
rect 33977 8412 34005 8443
rect 34164 8424 34192 8452
rect 34241 8449 34253 8483
rect 34287 8480 34299 8483
rect 34514 8480 34520 8492
rect 34287 8452 34520 8480
rect 34287 8449 34299 8452
rect 34241 8443 34299 8449
rect 34514 8440 34520 8452
rect 34572 8480 34578 8492
rect 35161 8483 35219 8489
rect 35161 8480 35173 8483
rect 34572 8452 35173 8480
rect 34572 8440 34578 8452
rect 35161 8449 35173 8452
rect 35207 8449 35219 8483
rect 35161 8443 35219 8449
rect 35250 8440 35256 8492
rect 35308 8480 35314 8492
rect 35434 8480 35440 8492
rect 35308 8452 35353 8480
rect 35395 8452 35440 8480
rect 35308 8440 35314 8452
rect 35434 8440 35440 8452
rect 35492 8440 35498 8492
rect 35618 8480 35624 8492
rect 35579 8452 35624 8480
rect 35618 8440 35624 8452
rect 35676 8440 35682 8492
rect 35894 8440 35900 8492
rect 35952 8480 35958 8492
rect 36464 8489 36492 8520
rect 36556 8520 37596 8548
rect 36556 8489 36584 8520
rect 42978 8508 42984 8560
rect 43036 8548 43042 8560
rect 45649 8551 45707 8557
rect 45649 8548 45661 8551
rect 43036 8520 45661 8548
rect 43036 8508 43042 8520
rect 45649 8517 45661 8520
rect 45695 8517 45707 8551
rect 46198 8548 46204 8560
rect 46159 8520 46204 8548
rect 45649 8511 45707 8517
rect 46198 8508 46204 8520
rect 46256 8508 46262 8560
rect 46566 8508 46572 8560
rect 46624 8548 46630 8560
rect 50246 8548 50252 8560
rect 46624 8520 50252 8548
rect 46624 8508 46630 8520
rect 36357 8483 36415 8489
rect 36357 8480 36369 8483
rect 35952 8452 36369 8480
rect 35952 8440 35958 8452
rect 36357 8449 36369 8452
rect 36403 8449 36415 8483
rect 36357 8443 36415 8449
rect 36449 8483 36507 8489
rect 36449 8449 36461 8483
rect 36495 8449 36507 8483
rect 36449 8443 36507 8449
rect 36541 8483 36599 8489
rect 36541 8449 36553 8483
rect 36587 8449 36599 8483
rect 36722 8480 36728 8492
rect 36683 8452 36728 8480
rect 36541 8443 36599 8449
rect 36722 8440 36728 8452
rect 36780 8440 36786 8492
rect 37734 8480 37740 8492
rect 37695 8452 37740 8480
rect 37734 8440 37740 8452
rect 37792 8440 37798 8492
rect 37921 8483 37979 8489
rect 37921 8449 37933 8483
rect 37967 8480 37979 8483
rect 38194 8480 38200 8492
rect 37967 8452 38200 8480
rect 37967 8449 37979 8452
rect 37921 8443 37979 8449
rect 38194 8440 38200 8452
rect 38252 8440 38258 8492
rect 38562 8440 38568 8492
rect 38620 8480 38626 8492
rect 38749 8483 38807 8489
rect 38749 8480 38761 8483
rect 38620 8452 38761 8480
rect 38620 8440 38626 8452
rect 38749 8449 38761 8452
rect 38795 8449 38807 8483
rect 39390 8480 39396 8492
rect 39351 8452 39396 8480
rect 38749 8443 38807 8449
rect 34146 8412 34152 8424
rect 33744 8384 34005 8412
rect 34059 8384 34152 8412
rect 33744 8372 33750 8384
rect 26418 8304 26424 8356
rect 26476 8344 26482 8356
rect 27525 8347 27583 8353
rect 27525 8344 27537 8347
rect 26476 8316 27537 8344
rect 26476 8304 26482 8316
rect 27525 8313 27537 8316
rect 27571 8344 27583 8347
rect 28350 8344 28356 8356
rect 27571 8316 28356 8344
rect 27571 8313 27583 8316
rect 27525 8307 27583 8313
rect 28350 8304 28356 8316
rect 28408 8304 28414 8356
rect 29089 8347 29147 8353
rect 29089 8313 29101 8347
rect 29135 8344 29147 8347
rect 29178 8344 29184 8356
rect 29135 8316 29184 8344
rect 29135 8313 29147 8316
rect 29089 8307 29147 8313
rect 29178 8304 29184 8316
rect 29236 8304 29242 8356
rect 30006 8304 30012 8356
rect 30064 8344 30070 8356
rect 34072 8344 34100 8384
rect 34146 8372 34152 8384
rect 34204 8372 34210 8424
rect 34698 8372 34704 8424
rect 34756 8412 34762 8424
rect 34977 8415 35035 8421
rect 34977 8412 34989 8415
rect 34756 8384 34989 8412
rect 34756 8372 34762 8384
rect 34977 8381 34989 8384
rect 35023 8381 35035 8415
rect 34977 8375 35035 8381
rect 37274 8372 37280 8424
rect 37332 8412 37338 8424
rect 38473 8415 38531 8421
rect 38473 8412 38485 8415
rect 37332 8384 38485 8412
rect 37332 8372 37338 8384
rect 38473 8381 38485 8384
rect 38519 8412 38531 8415
rect 38654 8412 38660 8424
rect 38519 8384 38660 8412
rect 38519 8381 38531 8384
rect 38473 8375 38531 8381
rect 38654 8372 38660 8384
rect 38712 8372 38718 8424
rect 38764 8412 38792 8443
rect 39390 8440 39396 8452
rect 39448 8440 39454 8492
rect 39574 8480 39580 8492
rect 39535 8452 39580 8480
rect 39574 8440 39580 8452
rect 39632 8440 39638 8492
rect 40586 8480 40592 8492
rect 40547 8452 40592 8480
rect 40586 8440 40592 8452
rect 40644 8440 40650 8492
rect 41417 8483 41475 8489
rect 41417 8449 41429 8483
rect 41463 8449 41475 8483
rect 41782 8480 41788 8492
rect 41743 8452 41788 8480
rect 41417 8443 41475 8449
rect 40313 8415 40371 8421
rect 40313 8412 40325 8415
rect 38764 8384 40325 8412
rect 40313 8381 40325 8384
rect 40359 8381 40371 8415
rect 41432 8412 41460 8443
rect 41782 8440 41788 8452
rect 41840 8440 41846 8492
rect 42061 8483 42119 8489
rect 42061 8449 42073 8483
rect 42107 8480 42119 8483
rect 42150 8480 42156 8492
rect 42107 8452 42156 8480
rect 42107 8449 42119 8452
rect 42061 8443 42119 8449
rect 42150 8440 42156 8452
rect 42208 8480 42214 8492
rect 42705 8483 42763 8489
rect 42705 8480 42717 8483
rect 42208 8452 42717 8480
rect 42208 8440 42214 8452
rect 42705 8449 42717 8452
rect 42751 8480 42763 8483
rect 42751 8452 43484 8480
rect 42751 8449 42763 8452
rect 42705 8443 42763 8449
rect 42978 8412 42984 8424
rect 41432 8384 42984 8412
rect 40313 8375 40371 8381
rect 42978 8372 42984 8384
rect 43036 8372 43042 8424
rect 43162 8412 43168 8424
rect 43123 8384 43168 8412
rect 43162 8372 43168 8384
rect 43220 8372 43226 8424
rect 43456 8412 43484 8452
rect 43530 8440 43536 8492
rect 43588 8480 43594 8492
rect 43588 8452 43633 8480
rect 43588 8440 43594 8452
rect 44082 8440 44088 8492
rect 44140 8480 44146 8492
rect 44361 8483 44419 8489
rect 44361 8480 44373 8483
rect 44140 8452 44373 8480
rect 44140 8440 44146 8452
rect 44361 8449 44373 8452
rect 44407 8449 44419 8483
rect 44361 8443 44419 8449
rect 44910 8440 44916 8492
rect 44968 8480 44974 8492
rect 45189 8483 45247 8489
rect 45189 8480 45201 8483
rect 44968 8452 45201 8480
rect 44968 8440 44974 8452
rect 45189 8449 45201 8452
rect 45235 8480 45247 8483
rect 45370 8480 45376 8492
rect 45235 8452 45376 8480
rect 45235 8449 45247 8452
rect 45189 8443 45247 8449
rect 45370 8440 45376 8452
rect 45428 8440 45434 8492
rect 45465 8483 45523 8489
rect 45465 8449 45477 8483
rect 45511 8449 45523 8483
rect 45465 8443 45523 8449
rect 44450 8412 44456 8424
rect 43456 8384 44312 8412
rect 44411 8384 44456 8412
rect 30064 8316 34100 8344
rect 30064 8304 30070 8316
rect 34606 8304 34612 8356
rect 34664 8344 34670 8356
rect 35345 8347 35403 8353
rect 35345 8344 35357 8347
rect 34664 8316 35357 8344
rect 34664 8304 34670 8316
rect 35345 8313 35357 8316
rect 35391 8313 35403 8347
rect 35345 8307 35403 8313
rect 35526 8304 35532 8356
rect 35584 8344 35590 8356
rect 39761 8347 39819 8353
rect 39761 8344 39773 8347
rect 35584 8316 39773 8344
rect 35584 8304 35590 8316
rect 39761 8313 39773 8316
rect 39807 8313 39819 8347
rect 40770 8344 40776 8356
rect 40731 8316 40776 8344
rect 39761 8307 39819 8313
rect 40770 8304 40776 8316
rect 40828 8304 40834 8356
rect 41509 8347 41567 8353
rect 41509 8313 41521 8347
rect 41555 8344 41567 8347
rect 41598 8344 41604 8356
rect 41555 8316 41604 8344
rect 41555 8313 41567 8316
rect 41509 8307 41567 8313
rect 41598 8304 41604 8316
rect 41656 8304 41662 8356
rect 44284 8344 44312 8384
rect 44450 8372 44456 8384
rect 44508 8372 44514 8424
rect 44542 8372 44548 8424
rect 44600 8412 44606 8424
rect 44600 8384 44645 8412
rect 44600 8372 44606 8384
rect 45480 8344 45508 8443
rect 46014 8440 46020 8492
rect 46072 8480 46078 8492
rect 46109 8483 46167 8489
rect 46109 8480 46121 8483
rect 46072 8452 46121 8480
rect 46072 8440 46078 8452
rect 46109 8449 46121 8452
rect 46155 8449 46167 8483
rect 46109 8443 46167 8449
rect 46293 8483 46351 8489
rect 46293 8449 46305 8483
rect 46339 8480 46351 8483
rect 46658 8480 46664 8492
rect 46339 8452 46664 8480
rect 46339 8449 46351 8452
rect 46293 8443 46351 8449
rect 46658 8440 46664 8452
rect 46716 8440 46722 8492
rect 46842 8440 46848 8492
rect 46900 8480 46906 8492
rect 47136 8489 47256 8490
rect 46937 8483 46995 8489
rect 46937 8480 46949 8483
rect 46900 8452 46949 8480
rect 46900 8440 46906 8452
rect 46937 8449 46949 8452
rect 46983 8449 46995 8483
rect 46937 8443 46995 8449
rect 47121 8483 47256 8489
rect 47121 8449 47133 8483
rect 47167 8480 47256 8483
rect 47578 8480 47584 8492
rect 47167 8462 47584 8480
rect 47167 8449 47179 8462
rect 47228 8452 47584 8462
rect 47121 8443 47179 8449
rect 45554 8372 45560 8424
rect 45612 8412 45618 8424
rect 46952 8412 46980 8443
rect 47578 8440 47584 8452
rect 47636 8440 47642 8492
rect 48041 8483 48099 8489
rect 48041 8449 48053 8483
rect 48087 8449 48099 8483
rect 48041 8443 48099 8449
rect 48056 8412 48084 8443
rect 48130 8440 48136 8492
rect 48188 8480 48194 8492
rect 49602 8480 49608 8492
rect 48188 8452 49608 8480
rect 48188 8440 48194 8452
rect 49602 8440 49608 8452
rect 49660 8440 49666 8492
rect 49712 8489 49740 8520
rect 50246 8508 50252 8520
rect 50304 8508 50310 8560
rect 51442 8508 51448 8560
rect 51500 8548 51506 8560
rect 51629 8551 51687 8557
rect 51629 8548 51641 8551
rect 51500 8520 51641 8548
rect 51500 8508 51506 8520
rect 51629 8517 51641 8520
rect 51675 8517 51687 8551
rect 51629 8511 51687 8517
rect 54570 8508 54576 8560
rect 54628 8548 54634 8560
rect 56965 8551 57023 8557
rect 56965 8548 56977 8551
rect 54628 8520 56977 8548
rect 54628 8508 54634 8520
rect 56965 8517 56977 8520
rect 57011 8517 57023 8551
rect 56965 8511 57023 8517
rect 49697 8483 49755 8489
rect 49697 8449 49709 8483
rect 49743 8449 49755 8483
rect 50062 8480 50068 8492
rect 50023 8452 50068 8480
rect 49697 8443 49755 8449
rect 50062 8440 50068 8452
rect 50120 8440 50126 8492
rect 51813 8483 51871 8489
rect 51813 8480 51825 8483
rect 51460 8452 51825 8480
rect 51460 8424 51488 8452
rect 51813 8449 51825 8452
rect 51859 8449 51871 8483
rect 51813 8443 51871 8449
rect 51997 8483 52055 8489
rect 51997 8449 52009 8483
rect 52043 8449 52055 8483
rect 51997 8443 52055 8449
rect 52089 8483 52147 8489
rect 52089 8449 52101 8483
rect 52135 8480 52147 8483
rect 52178 8480 52184 8492
rect 52135 8452 52184 8480
rect 52135 8449 52147 8452
rect 52089 8443 52147 8449
rect 48314 8412 48320 8424
rect 45612 8384 48084 8412
rect 48275 8384 48320 8412
rect 45612 8372 45618 8384
rect 48314 8372 48320 8384
rect 48372 8372 48378 8424
rect 49786 8412 49792 8424
rect 49747 8384 49792 8412
rect 49786 8372 49792 8384
rect 49844 8372 49850 8424
rect 49881 8415 49939 8421
rect 49881 8381 49893 8415
rect 49927 8412 49939 8415
rect 50154 8412 50160 8424
rect 49927 8384 50160 8412
rect 49927 8381 49939 8384
rect 49881 8375 49939 8381
rect 46566 8344 46572 8356
rect 44284 8316 46572 8344
rect 46566 8304 46572 8316
rect 46624 8304 46630 8356
rect 47118 8344 47124 8356
rect 47079 8316 47124 8344
rect 47118 8304 47124 8316
rect 47176 8304 47182 8356
rect 48225 8347 48283 8353
rect 48225 8313 48237 8347
rect 48271 8344 48283 8347
rect 49421 8347 49479 8353
rect 49421 8344 49433 8347
rect 48271 8316 49433 8344
rect 48271 8313 48283 8316
rect 48225 8307 48283 8313
rect 49421 8313 49433 8316
rect 49467 8313 49479 8347
rect 49421 8307 49479 8313
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 26878 8276 26884 8288
rect 2372 8248 26884 8276
rect 2372 8236 2378 8248
rect 26878 8236 26884 8248
rect 26936 8236 26942 8288
rect 29270 8236 29276 8288
rect 29328 8276 29334 8288
rect 29914 8276 29920 8288
rect 29328 8248 29920 8276
rect 29328 8236 29334 8248
rect 29914 8236 29920 8248
rect 29972 8236 29978 8288
rect 33594 8276 33600 8288
rect 33555 8248 33600 8276
rect 33594 8236 33600 8248
rect 33652 8236 33658 8288
rect 36081 8279 36139 8285
rect 36081 8245 36093 8279
rect 36127 8276 36139 8279
rect 36170 8276 36176 8288
rect 36127 8248 36176 8276
rect 36127 8245 36139 8248
rect 36081 8239 36139 8245
rect 36170 8236 36176 8248
rect 36228 8236 36234 8288
rect 37366 8236 37372 8288
rect 37424 8276 37430 8288
rect 38565 8279 38623 8285
rect 38565 8276 38577 8279
rect 37424 8248 38577 8276
rect 37424 8236 37430 8248
rect 38565 8245 38577 8248
rect 38611 8276 38623 8279
rect 38838 8276 38844 8288
rect 38611 8248 38844 8276
rect 38611 8245 38623 8248
rect 38565 8239 38623 8245
rect 38838 8236 38844 8248
rect 38896 8236 38902 8288
rect 40402 8276 40408 8288
rect 40363 8248 40408 8276
rect 40402 8236 40408 8248
rect 40460 8236 40466 8288
rect 45278 8276 45284 8288
rect 45239 8248 45284 8276
rect 45278 8236 45284 8248
rect 45336 8236 45342 8288
rect 46934 8236 46940 8288
rect 46992 8276 46998 8288
rect 48130 8276 48136 8288
rect 46992 8248 48136 8276
rect 46992 8236 46998 8248
rect 48130 8236 48136 8248
rect 48188 8236 48194 8288
rect 49694 8236 49700 8288
rect 49752 8276 49758 8288
rect 49988 8276 50016 8384
rect 50154 8372 50160 8384
rect 50212 8372 50218 8424
rect 50525 8415 50583 8421
rect 50525 8381 50537 8415
rect 50571 8381 50583 8415
rect 50525 8375 50583 8381
rect 50540 8344 50568 8375
rect 50798 8372 50804 8424
rect 50856 8412 50862 8424
rect 50893 8415 50951 8421
rect 50893 8412 50905 8415
rect 50856 8384 50905 8412
rect 50856 8372 50862 8384
rect 50893 8381 50905 8384
rect 50939 8381 50951 8415
rect 50893 8375 50951 8381
rect 51442 8372 51448 8424
rect 51500 8372 51506 8424
rect 51534 8372 51540 8424
rect 51592 8412 51598 8424
rect 51902 8412 51908 8424
rect 51592 8384 51908 8412
rect 51592 8372 51598 8384
rect 51902 8372 51908 8384
rect 51960 8412 51966 8424
rect 52012 8412 52040 8443
rect 52178 8440 52184 8452
rect 52236 8440 52242 8492
rect 52914 8480 52920 8492
rect 52875 8452 52920 8480
rect 52914 8440 52920 8452
rect 52972 8440 52978 8492
rect 53377 8483 53435 8489
rect 53377 8449 53389 8483
rect 53423 8449 53435 8483
rect 54665 8483 54723 8489
rect 54665 8480 54677 8483
rect 53377 8443 53435 8449
rect 53484 8452 54677 8480
rect 51960 8384 52040 8412
rect 52196 8412 52224 8440
rect 53392 8412 53420 8443
rect 52196 8384 53420 8412
rect 51960 8372 51966 8384
rect 50614 8344 50620 8356
rect 50527 8316 50620 8344
rect 50614 8304 50620 8316
rect 50672 8344 50678 8356
rect 53484 8344 53512 8452
rect 54665 8449 54677 8452
rect 54711 8480 54723 8483
rect 54846 8480 54852 8492
rect 54711 8452 54852 8480
rect 54711 8449 54723 8452
rect 54665 8443 54723 8449
rect 54846 8440 54852 8452
rect 54904 8480 54910 8492
rect 55309 8483 55367 8489
rect 55309 8480 55321 8483
rect 54904 8452 55321 8480
rect 54904 8440 54910 8452
rect 55309 8449 55321 8452
rect 55355 8449 55367 8483
rect 55309 8443 55367 8449
rect 55401 8483 55459 8489
rect 55401 8449 55413 8483
rect 55447 8480 55459 8483
rect 55490 8480 55496 8492
rect 55447 8452 55496 8480
rect 55447 8449 55459 8452
rect 55401 8443 55459 8449
rect 53653 8415 53711 8421
rect 53653 8381 53665 8415
rect 53699 8412 53711 8415
rect 54018 8412 54024 8424
rect 53699 8384 54024 8412
rect 53699 8381 53711 8384
rect 53653 8375 53711 8381
rect 54018 8372 54024 8384
rect 54076 8372 54082 8424
rect 55416 8412 55444 8443
rect 55490 8440 55496 8452
rect 55548 8440 55554 8492
rect 55769 8483 55827 8489
rect 55769 8449 55781 8483
rect 55815 8480 55827 8483
rect 56042 8480 56048 8492
rect 55815 8452 56048 8480
rect 55815 8449 55827 8452
rect 55769 8443 55827 8449
rect 56042 8440 56048 8452
rect 56100 8440 56106 8492
rect 56410 8480 56416 8492
rect 56371 8452 56416 8480
rect 56410 8440 56416 8452
rect 56468 8480 56474 8492
rect 57146 8480 57152 8492
rect 56468 8452 57152 8480
rect 56468 8440 56474 8452
rect 57146 8440 57152 8452
rect 57204 8440 57210 8492
rect 54312 8384 55444 8412
rect 54312 8356 54340 8384
rect 50672 8316 53512 8344
rect 54205 8347 54263 8353
rect 50672 8304 50678 8316
rect 54205 8313 54217 8347
rect 54251 8344 54263 8347
rect 54294 8344 54300 8356
rect 54251 8316 54300 8344
rect 54251 8313 54263 8316
rect 54205 8307 54263 8313
rect 54294 8304 54300 8316
rect 54352 8304 54358 8356
rect 55398 8344 55404 8356
rect 55359 8316 55404 8344
rect 55398 8304 55404 8316
rect 55456 8304 55462 8356
rect 50890 8276 50896 8288
rect 49752 8248 50016 8276
rect 50851 8248 50896 8276
rect 49752 8236 49758 8248
rect 50890 8236 50896 8248
rect 50948 8236 50954 8288
rect 50982 8236 50988 8288
rect 51040 8276 51046 8288
rect 54386 8276 54392 8288
rect 51040 8248 54392 8276
rect 51040 8236 51046 8248
rect 54386 8236 54392 8248
rect 54444 8236 54450 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 24581 8075 24639 8081
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 25314 8072 25320 8084
rect 24627 8044 25320 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 25314 8032 25320 8044
rect 25372 8032 25378 8084
rect 27430 8072 27436 8084
rect 27391 8044 27436 8072
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 27798 8032 27804 8084
rect 27856 8072 27862 8084
rect 29917 8075 29975 8081
rect 29917 8072 29929 8075
rect 27856 8044 29929 8072
rect 27856 8032 27862 8044
rect 29917 8041 29929 8044
rect 29963 8072 29975 8075
rect 32950 8072 32956 8084
rect 29963 8044 32956 8072
rect 29963 8041 29975 8044
rect 29917 8035 29975 8041
rect 32950 8032 32956 8044
rect 33008 8032 33014 8084
rect 33229 8075 33287 8081
rect 33229 8041 33241 8075
rect 33275 8072 33287 8075
rect 33686 8072 33692 8084
rect 33275 8044 33692 8072
rect 33275 8041 33287 8044
rect 33229 8035 33287 8041
rect 33686 8032 33692 8044
rect 33744 8072 33750 8084
rect 34606 8072 34612 8084
rect 33744 8044 34612 8072
rect 33744 8032 33750 8044
rect 34606 8032 34612 8044
rect 34664 8032 34670 8084
rect 35253 8075 35311 8081
rect 35253 8041 35265 8075
rect 35299 8072 35311 8075
rect 35434 8072 35440 8084
rect 35299 8044 35440 8072
rect 35299 8041 35311 8044
rect 35253 8035 35311 8041
rect 35434 8032 35440 8044
rect 35492 8032 35498 8084
rect 35618 8032 35624 8084
rect 35676 8072 35682 8084
rect 35805 8075 35863 8081
rect 35805 8072 35817 8075
rect 35676 8044 35817 8072
rect 35676 8032 35682 8044
rect 35805 8041 35817 8044
rect 35851 8041 35863 8075
rect 35986 8072 35992 8084
rect 35947 8044 35992 8072
rect 35805 8035 35863 8041
rect 35986 8032 35992 8044
rect 36044 8032 36050 8084
rect 36262 8032 36268 8084
rect 36320 8072 36326 8084
rect 36817 8075 36875 8081
rect 36817 8072 36829 8075
rect 36320 8044 36829 8072
rect 36320 8032 36326 8044
rect 36817 8041 36829 8044
rect 36863 8072 36875 8075
rect 37734 8072 37740 8084
rect 36863 8044 37740 8072
rect 36863 8041 36875 8044
rect 36817 8035 36875 8041
rect 37734 8032 37740 8044
rect 37792 8032 37798 8084
rect 38654 8032 38660 8084
rect 38712 8072 38718 8084
rect 38749 8075 38807 8081
rect 38749 8072 38761 8075
rect 38712 8044 38761 8072
rect 38712 8032 38718 8044
rect 38749 8041 38761 8044
rect 38795 8072 38807 8075
rect 39022 8072 39028 8084
rect 38795 8044 39028 8072
rect 38795 8041 38807 8044
rect 38749 8035 38807 8041
rect 39022 8032 39028 8044
rect 39080 8032 39086 8084
rect 40405 8075 40463 8081
rect 40405 8041 40417 8075
rect 40451 8072 40463 8075
rect 40494 8072 40500 8084
rect 40451 8044 40500 8072
rect 40451 8041 40463 8044
rect 40405 8035 40463 8041
rect 40494 8032 40500 8044
rect 40552 8032 40558 8084
rect 40954 8072 40960 8084
rect 40915 8044 40960 8072
rect 40954 8032 40960 8044
rect 41012 8032 41018 8084
rect 41322 8032 41328 8084
rect 41380 8072 41386 8084
rect 42061 8075 42119 8081
rect 42061 8072 42073 8075
rect 41380 8044 42073 8072
rect 41380 8032 41386 8044
rect 42061 8041 42073 8044
rect 42107 8072 42119 8075
rect 42518 8072 42524 8084
rect 42107 8044 42524 8072
rect 42107 8041 42119 8044
rect 42061 8035 42119 8041
rect 42518 8032 42524 8044
rect 42576 8032 42582 8084
rect 45833 8075 45891 8081
rect 45833 8041 45845 8075
rect 45879 8072 45891 8075
rect 46474 8072 46480 8084
rect 45879 8044 46480 8072
rect 45879 8041 45891 8044
rect 45833 8035 45891 8041
rect 46474 8032 46480 8044
rect 46532 8032 46538 8084
rect 46566 8032 46572 8084
rect 46624 8072 46630 8084
rect 47854 8072 47860 8084
rect 46624 8044 47860 8072
rect 46624 8032 46630 8044
rect 47854 8032 47860 8044
rect 47912 8032 47918 8084
rect 48317 8075 48375 8081
rect 48317 8041 48329 8075
rect 48363 8072 48375 8075
rect 48406 8072 48412 8084
rect 48363 8044 48412 8072
rect 48363 8041 48375 8044
rect 48317 8035 48375 8041
rect 48406 8032 48412 8044
rect 48464 8032 48470 8084
rect 49789 8075 49847 8081
rect 49789 8041 49801 8075
rect 49835 8072 49847 8075
rect 49878 8072 49884 8084
rect 49835 8044 49884 8072
rect 49835 8041 49847 8044
rect 49789 8035 49847 8041
rect 49878 8032 49884 8044
rect 49936 8032 49942 8084
rect 50798 8032 50804 8084
rect 50856 8072 50862 8084
rect 51810 8072 51816 8084
rect 50856 8044 51672 8072
rect 51771 8044 51816 8072
rect 50856 8032 50862 8044
rect 25774 8004 25780 8016
rect 25735 7976 25780 8004
rect 25774 7964 25780 7976
rect 25832 7964 25838 8016
rect 27065 8007 27123 8013
rect 27065 8004 27077 8007
rect 26160 7976 27077 8004
rect 25501 7939 25559 7945
rect 25501 7905 25513 7939
rect 25547 7936 25559 7939
rect 26160 7936 26188 7976
rect 27065 7973 27077 7976
rect 27111 8004 27123 8007
rect 27246 8004 27252 8016
rect 27111 7976 27252 8004
rect 27111 7973 27123 7976
rect 27065 7967 27123 7973
rect 27246 7964 27252 7976
rect 27304 7964 27310 8016
rect 28810 7964 28816 8016
rect 28868 8004 28874 8016
rect 32766 8004 32772 8016
rect 28868 7976 32772 8004
rect 28868 7964 28874 7976
rect 32766 7964 32772 7976
rect 32824 7964 32830 8016
rect 33134 7964 33140 8016
rect 33192 8004 33198 8016
rect 33781 8007 33839 8013
rect 33781 8004 33793 8007
rect 33192 7976 33793 8004
rect 33192 7964 33198 7976
rect 33781 7973 33793 7976
rect 33827 7973 33839 8007
rect 38930 8004 38936 8016
rect 33781 7967 33839 7973
rect 33888 7976 38654 8004
rect 38843 7976 38936 8004
rect 26510 7936 26516 7948
rect 25547 7908 26188 7936
rect 26252 7908 26516 7936
rect 25547 7905 25559 7908
rect 25501 7899 25559 7905
rect 25222 7828 25228 7880
rect 25280 7868 25286 7880
rect 25406 7877 25412 7880
rect 25384 7871 25412 7877
rect 25280 7840 25325 7868
rect 25280 7828 25286 7840
rect 25384 7837 25396 7871
rect 25384 7831 25412 7837
rect 25406 7828 25412 7831
rect 25464 7828 25470 7880
rect 26252 7877 26280 7908
rect 26510 7896 26516 7908
rect 26568 7936 26574 7948
rect 26786 7936 26792 7948
rect 26568 7908 26792 7936
rect 26568 7896 26574 7908
rect 26786 7896 26792 7908
rect 26844 7896 26850 7948
rect 26878 7896 26884 7948
rect 26936 7936 26942 7948
rect 33888 7936 33916 7976
rect 35158 7936 35164 7948
rect 26936 7908 33916 7936
rect 34992 7908 35164 7936
rect 26936 7896 26942 7908
rect 26237 7871 26295 7877
rect 26237 7837 26249 7871
rect 26283 7837 26295 7871
rect 26237 7831 26295 7837
rect 26421 7871 26479 7877
rect 26421 7837 26433 7871
rect 26467 7837 26479 7871
rect 26970 7868 26976 7880
rect 26931 7840 26976 7868
rect 26421 7831 26479 7837
rect 26436 7732 26464 7831
rect 26970 7828 26976 7840
rect 27028 7828 27034 7880
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7837 27307 7871
rect 27249 7831 27307 7837
rect 27985 7871 28043 7877
rect 27985 7837 27997 7871
rect 28031 7868 28043 7871
rect 28534 7868 28540 7880
rect 28031 7840 28540 7868
rect 28031 7837 28043 7840
rect 27985 7831 28043 7837
rect 27264 7800 27292 7831
rect 28534 7828 28540 7840
rect 28592 7828 28598 7880
rect 28813 7871 28871 7877
rect 28813 7837 28825 7871
rect 28859 7868 28871 7871
rect 29086 7868 29092 7880
rect 28859 7840 29092 7868
rect 28859 7837 28871 7840
rect 28813 7831 28871 7837
rect 29086 7828 29092 7840
rect 29144 7828 29150 7880
rect 29546 7828 29552 7880
rect 29604 7868 29610 7880
rect 29733 7871 29791 7877
rect 29733 7868 29745 7871
rect 29604 7840 29745 7868
rect 29604 7828 29610 7840
rect 29733 7837 29745 7840
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 29822 7828 29828 7880
rect 29880 7868 29886 7880
rect 31389 7871 31447 7877
rect 29880 7840 29925 7868
rect 29880 7828 29886 7840
rect 31389 7837 31401 7871
rect 31435 7870 31447 7871
rect 31478 7870 31484 7880
rect 31435 7842 31484 7870
rect 31435 7837 31447 7842
rect 31389 7831 31447 7837
rect 31478 7828 31484 7842
rect 31536 7828 31542 7880
rect 31754 7868 31760 7880
rect 31715 7840 31760 7868
rect 31754 7828 31760 7840
rect 31812 7828 31818 7880
rect 32122 7868 32128 7880
rect 32083 7840 32128 7868
rect 32122 7828 32128 7840
rect 32180 7828 32186 7880
rect 32490 7828 32496 7880
rect 32548 7868 32554 7880
rect 33134 7868 33140 7880
rect 32548 7840 33140 7868
rect 32548 7828 32554 7840
rect 33134 7828 33140 7840
rect 33192 7828 33198 7880
rect 33229 7871 33287 7877
rect 33229 7837 33241 7871
rect 33275 7837 33287 7871
rect 33229 7831 33287 7837
rect 27522 7800 27528 7812
rect 27264 7772 27528 7800
rect 27522 7760 27528 7772
rect 27580 7800 27586 7812
rect 28445 7803 28503 7809
rect 28445 7800 28457 7803
rect 27580 7772 28457 7800
rect 27580 7760 27586 7772
rect 28445 7769 28457 7772
rect 28491 7800 28503 7803
rect 28902 7800 28908 7812
rect 28491 7772 28908 7800
rect 28491 7769 28503 7772
rect 28445 7763 28503 7769
rect 28902 7760 28908 7772
rect 28960 7760 28966 7812
rect 30282 7760 30288 7812
rect 30340 7800 30346 7812
rect 30340 7772 31432 7800
rect 30340 7760 30346 7772
rect 28258 7732 28264 7744
rect 26436 7704 28264 7732
rect 28258 7692 28264 7704
rect 28316 7692 28322 7744
rect 28994 7692 29000 7744
rect 29052 7732 29058 7744
rect 29822 7732 29828 7744
rect 29052 7704 29828 7732
rect 29052 7692 29058 7704
rect 29822 7692 29828 7704
rect 29880 7692 29886 7744
rect 30101 7735 30159 7741
rect 30101 7701 30113 7735
rect 30147 7732 30159 7735
rect 30466 7732 30472 7744
rect 30147 7704 30472 7732
rect 30147 7701 30159 7704
rect 30101 7695 30159 7701
rect 30466 7692 30472 7704
rect 30524 7692 30530 7744
rect 30650 7732 30656 7744
rect 30611 7704 30656 7732
rect 30650 7692 30656 7704
rect 30708 7692 30714 7744
rect 31110 7692 31116 7744
rect 31168 7732 31174 7744
rect 31297 7735 31355 7741
rect 31297 7732 31309 7735
rect 31168 7704 31309 7732
rect 31168 7692 31174 7704
rect 31297 7701 31309 7704
rect 31343 7701 31355 7735
rect 31404 7732 31432 7772
rect 32306 7760 32312 7812
rect 32364 7800 32370 7812
rect 33244 7800 33272 7831
rect 33594 7828 33600 7880
rect 33652 7868 33658 7880
rect 33781 7871 33839 7877
rect 33781 7868 33793 7871
rect 33652 7840 33793 7868
rect 33652 7828 33658 7840
rect 33781 7837 33793 7840
rect 33827 7837 33839 7871
rect 34054 7868 34060 7880
rect 34015 7840 34060 7868
rect 33781 7831 33839 7837
rect 34054 7828 34060 7840
rect 34112 7828 34118 7880
rect 34992 7800 35020 7908
rect 35158 7896 35164 7908
rect 35216 7896 35222 7948
rect 35345 7939 35403 7945
rect 35345 7905 35357 7939
rect 35391 7936 35403 7939
rect 35391 7908 36216 7936
rect 35391 7905 35403 7908
rect 35345 7899 35403 7905
rect 36188 7880 36216 7908
rect 35069 7871 35127 7877
rect 35069 7837 35081 7871
rect 35115 7837 35127 7871
rect 35069 7831 35127 7837
rect 32364 7772 35020 7800
rect 35084 7800 35112 7831
rect 35894 7828 35900 7880
rect 35952 7868 35958 7880
rect 35989 7871 36047 7877
rect 35989 7868 36001 7871
rect 35952 7840 36001 7868
rect 35952 7828 35958 7840
rect 35989 7837 36001 7840
rect 36035 7837 36047 7871
rect 36170 7868 36176 7880
rect 36131 7840 36176 7868
rect 35989 7831 36047 7837
rect 36170 7828 36176 7840
rect 36228 7828 36234 7880
rect 36722 7868 36728 7880
rect 36683 7840 36728 7868
rect 36722 7828 36728 7840
rect 36780 7828 36786 7880
rect 37642 7828 37648 7880
rect 37700 7868 37706 7880
rect 37737 7871 37795 7877
rect 37737 7868 37749 7871
rect 37700 7840 37749 7868
rect 37700 7828 37706 7840
rect 37737 7837 37749 7840
rect 37783 7837 37795 7871
rect 38010 7868 38016 7880
rect 37971 7840 38016 7868
rect 37737 7831 37795 7837
rect 38010 7828 38016 7840
rect 38068 7828 38074 7880
rect 38626 7868 38654 7976
rect 38930 7964 38936 7976
rect 38988 8004 38994 8016
rect 39390 8004 39396 8016
rect 38988 7976 39396 8004
rect 38988 7964 38994 7976
rect 39390 7964 39396 7976
rect 39448 7964 39454 8016
rect 40218 7964 40224 8016
rect 40276 8004 40282 8016
rect 41340 8004 41368 8032
rect 42794 8004 42800 8016
rect 40276 7976 41368 8004
rect 42755 7976 42800 8004
rect 40276 7964 40282 7976
rect 42794 7964 42800 7976
rect 42852 7964 42858 8016
rect 46382 7964 46388 8016
rect 46440 8004 46446 8016
rect 51166 8004 51172 8016
rect 46440 7976 51172 8004
rect 46440 7964 46446 7976
rect 51166 7964 51172 7976
rect 51224 7964 51230 8016
rect 51350 7964 51356 8016
rect 51408 7964 51414 8016
rect 51644 8004 51672 8044
rect 51810 8032 51816 8044
rect 51868 8032 51874 8084
rect 52086 8032 52092 8084
rect 52144 8072 52150 8084
rect 52641 8075 52699 8081
rect 52641 8072 52653 8075
rect 52144 8044 52653 8072
rect 52144 8032 52150 8044
rect 52641 8041 52653 8044
rect 52687 8041 52699 8075
rect 56042 8072 56048 8084
rect 52641 8035 52699 8041
rect 54588 8044 56048 8072
rect 51644 7976 52224 8004
rect 39209 7939 39267 7945
rect 39209 7905 39221 7939
rect 39255 7936 39267 7939
rect 39574 7936 39580 7948
rect 39255 7908 39580 7936
rect 39255 7905 39267 7908
rect 39209 7899 39267 7905
rect 39574 7896 39580 7908
rect 39632 7896 39638 7948
rect 42150 7936 42156 7948
rect 40144 7908 42156 7936
rect 40144 7877 40172 7908
rect 42150 7896 42156 7908
rect 42208 7896 42214 7948
rect 42702 7896 42708 7948
rect 42760 7936 42766 7948
rect 44082 7936 44088 7948
rect 42760 7908 44088 7936
rect 42760 7896 42766 7908
rect 40129 7871 40187 7877
rect 40129 7868 40141 7871
rect 38626 7840 40141 7868
rect 40129 7837 40141 7840
rect 40175 7837 40187 7871
rect 40129 7831 40187 7837
rect 41414 7828 41420 7880
rect 41472 7868 41478 7880
rect 42812 7877 42840 7908
rect 44082 7896 44088 7908
rect 44140 7896 44146 7948
rect 46750 7896 46756 7948
rect 46808 7936 46814 7948
rect 46808 7908 46888 7936
rect 46808 7896 46814 7908
rect 42613 7871 42671 7877
rect 42613 7868 42625 7871
rect 41472 7840 42625 7868
rect 41472 7828 41478 7840
rect 42613 7837 42625 7840
rect 42659 7837 42671 7871
rect 42613 7831 42671 7837
rect 42797 7871 42855 7877
rect 42797 7837 42809 7871
rect 42843 7837 42855 7871
rect 44266 7868 44272 7880
rect 42797 7831 42855 7837
rect 43732 7840 44272 7868
rect 36538 7800 36544 7812
rect 35084 7772 36544 7800
rect 32364 7760 32370 7772
rect 36538 7760 36544 7772
rect 36596 7760 36602 7812
rect 41598 7760 41604 7812
rect 41656 7800 41662 7812
rect 42812 7800 42840 7831
rect 41656 7772 42840 7800
rect 41656 7760 41662 7772
rect 33965 7735 34023 7741
rect 33965 7732 33977 7735
rect 31404 7704 33977 7732
rect 31297 7695 31355 7701
rect 33965 7701 33977 7704
rect 34011 7701 34023 7735
rect 38194 7732 38200 7744
rect 38155 7704 38200 7732
rect 33965 7695 34023 7701
rect 38194 7692 38200 7704
rect 38252 7692 38258 7744
rect 41506 7732 41512 7744
rect 41467 7704 41512 7732
rect 41506 7692 41512 7704
rect 41564 7692 41570 7744
rect 43254 7692 43260 7744
rect 43312 7732 43318 7744
rect 43732 7732 43760 7840
rect 44266 7828 44272 7840
rect 44324 7828 44330 7880
rect 44450 7828 44456 7880
rect 44508 7868 44514 7880
rect 46566 7868 46572 7880
rect 44508 7840 46572 7868
rect 44508 7828 44514 7840
rect 46566 7828 46572 7840
rect 46624 7828 46630 7880
rect 46860 7877 46888 7908
rect 47578 7896 47584 7948
rect 47636 7936 47642 7948
rect 49421 7939 49479 7945
rect 47636 7908 48314 7936
rect 47636 7896 47642 7908
rect 46661 7871 46719 7877
rect 46661 7837 46673 7871
rect 46707 7868 46719 7871
rect 46857 7871 46915 7877
rect 46707 7840 46796 7868
rect 46707 7837 46719 7840
rect 46661 7831 46719 7837
rect 43809 7803 43867 7809
rect 43809 7769 43821 7803
rect 43855 7800 43867 7803
rect 44542 7800 44548 7812
rect 43855 7772 44548 7800
rect 43855 7769 43867 7772
rect 43809 7763 43867 7769
rect 44542 7760 44548 7772
rect 44600 7760 44606 7812
rect 43901 7735 43959 7741
rect 43901 7732 43913 7735
rect 43312 7704 43913 7732
rect 43312 7692 43318 7704
rect 43901 7701 43913 7704
rect 43947 7701 43959 7735
rect 43901 7695 43959 7701
rect 44082 7692 44088 7744
rect 44140 7732 44146 7744
rect 45281 7735 45339 7741
rect 45281 7732 45293 7735
rect 44140 7704 45293 7732
rect 44140 7692 44146 7704
rect 45281 7701 45293 7704
rect 45327 7732 45339 7735
rect 45830 7732 45836 7744
rect 45327 7704 45836 7732
rect 45327 7701 45339 7704
rect 45281 7695 45339 7701
rect 45830 7692 45836 7704
rect 45888 7692 45894 7744
rect 46290 7692 46296 7744
rect 46348 7732 46354 7744
rect 46385 7735 46443 7741
rect 46385 7732 46397 7735
rect 46348 7704 46397 7732
rect 46348 7692 46354 7704
rect 46385 7701 46397 7704
rect 46431 7701 46443 7735
rect 46385 7695 46443 7701
rect 46474 7692 46480 7744
rect 46532 7732 46538 7744
rect 46768 7732 46796 7840
rect 46857 7837 46869 7871
rect 46903 7837 46915 7871
rect 46857 7831 46915 7837
rect 46947 7871 47005 7877
rect 46947 7837 46959 7871
rect 46993 7868 47005 7871
rect 47670 7868 47676 7880
rect 46993 7840 47676 7868
rect 46993 7837 47005 7840
rect 46947 7831 47005 7837
rect 47670 7828 47676 7840
rect 47728 7828 47734 7880
rect 47854 7868 47860 7880
rect 47815 7840 47860 7868
rect 47854 7828 47860 7840
rect 47912 7828 47918 7880
rect 47949 7871 48007 7877
rect 47949 7837 47961 7871
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 48041 7871 48099 7877
rect 48041 7837 48053 7871
rect 48087 7868 48099 7871
rect 48130 7868 48136 7880
rect 48087 7840 48136 7868
rect 48087 7837 48099 7840
rect 48041 7831 48099 7837
rect 46532 7704 46796 7732
rect 47688 7732 47716 7828
rect 47964 7800 47992 7831
rect 48130 7828 48136 7840
rect 48188 7828 48194 7880
rect 48286 7868 48314 7908
rect 49421 7905 49433 7939
rect 49467 7936 49479 7939
rect 49786 7936 49792 7948
rect 49467 7908 49792 7936
rect 49467 7905 49479 7908
rect 49421 7899 49479 7905
rect 49786 7896 49792 7908
rect 49844 7936 49850 7948
rect 50062 7936 50068 7948
rect 49844 7908 50068 7936
rect 49844 7896 49850 7908
rect 50062 7896 50068 7908
rect 50120 7896 50126 7948
rect 50709 7939 50767 7945
rect 50709 7905 50721 7939
rect 50755 7936 50767 7939
rect 50982 7936 50988 7948
rect 50755 7908 50988 7936
rect 50755 7905 50767 7908
rect 50709 7899 50767 7905
rect 50982 7896 50988 7908
rect 51040 7896 51046 7948
rect 51368 7936 51396 7964
rect 51902 7936 51908 7948
rect 51368 7908 51908 7936
rect 49326 7868 49332 7880
rect 48286 7840 49332 7868
rect 49326 7828 49332 7840
rect 49384 7828 49390 7880
rect 49510 7868 49516 7880
rect 49471 7840 49516 7868
rect 49510 7828 49516 7840
rect 49568 7828 49574 7880
rect 51368 7877 51396 7908
rect 51902 7896 51908 7908
rect 51960 7896 51966 7948
rect 49605 7871 49663 7877
rect 49605 7837 49617 7871
rect 49651 7868 49663 7871
rect 51261 7871 51319 7877
rect 49651 7840 49740 7868
rect 49651 7837 49663 7840
rect 49605 7831 49663 7837
rect 48222 7800 48228 7812
rect 47964 7772 48228 7800
rect 48222 7760 48228 7772
rect 48280 7760 48286 7812
rect 49712 7732 49740 7840
rect 51261 7837 51273 7871
rect 51307 7837 51319 7871
rect 51261 7831 51319 7837
rect 51353 7871 51411 7877
rect 51353 7837 51365 7871
rect 51399 7837 51411 7871
rect 51534 7868 51540 7880
rect 51495 7840 51540 7868
rect 51353 7831 51411 7837
rect 49878 7760 49884 7812
rect 49936 7800 49942 7812
rect 50433 7803 50491 7809
rect 50433 7800 50445 7803
rect 49936 7772 50445 7800
rect 49936 7760 49942 7772
rect 50433 7769 50445 7772
rect 50479 7769 50491 7803
rect 51276 7800 51304 7831
rect 51534 7828 51540 7840
rect 51592 7828 51598 7880
rect 51629 7871 51687 7877
rect 51629 7837 51641 7871
rect 51675 7868 51687 7871
rect 51994 7868 52000 7880
rect 51675 7840 52000 7868
rect 51675 7837 51687 7840
rect 51629 7831 51687 7837
rect 51994 7828 52000 7840
rect 52052 7828 52058 7880
rect 51442 7800 51448 7812
rect 51276 7772 51448 7800
rect 50433 7763 50491 7769
rect 51442 7760 51448 7772
rect 51500 7760 51506 7812
rect 52196 7800 52224 7976
rect 52270 7964 52276 8016
rect 52328 8004 52334 8016
rect 53561 8007 53619 8013
rect 53561 8004 53573 8007
rect 52328 7976 53573 8004
rect 52328 7964 52334 7976
rect 53561 7973 53573 7976
rect 53607 7973 53619 8007
rect 53561 7967 53619 7973
rect 53466 7936 53472 7948
rect 52840 7908 53472 7936
rect 52840 7877 52868 7908
rect 53466 7896 53472 7908
rect 53524 7896 53530 7948
rect 52825 7871 52883 7877
rect 52825 7837 52837 7871
rect 52871 7837 52883 7871
rect 53006 7868 53012 7880
rect 52967 7840 53012 7868
rect 52825 7831 52883 7837
rect 53006 7828 53012 7840
rect 53064 7828 53070 7880
rect 53101 7871 53159 7877
rect 53101 7837 53113 7871
rect 53147 7868 53159 7871
rect 53282 7868 53288 7880
rect 53147 7840 53288 7868
rect 53147 7837 53159 7840
rect 53101 7831 53159 7837
rect 53282 7828 53288 7840
rect 53340 7828 53346 7880
rect 53745 7871 53803 7877
rect 53745 7837 53757 7871
rect 53791 7837 53803 7871
rect 53745 7831 53803 7837
rect 53929 7871 53987 7877
rect 53929 7837 53941 7871
rect 53975 7868 53987 7871
rect 54110 7868 54116 7880
rect 53975 7840 54116 7868
rect 53975 7837 53987 7840
rect 53929 7831 53987 7837
rect 53650 7800 53656 7812
rect 52196 7772 53656 7800
rect 53650 7760 53656 7772
rect 53708 7760 53714 7812
rect 53760 7800 53788 7831
rect 54110 7828 54116 7840
rect 54168 7828 54174 7880
rect 54386 7868 54392 7880
rect 54347 7840 54392 7868
rect 54386 7828 54392 7840
rect 54444 7828 54450 7880
rect 54588 7877 54616 8044
rect 56042 8032 56048 8044
rect 56100 8072 56106 8084
rect 56137 8075 56195 8081
rect 56137 8072 56149 8075
rect 56100 8044 56149 8072
rect 56100 8032 56106 8044
rect 56137 8041 56149 8044
rect 56183 8041 56195 8075
rect 57422 8072 57428 8084
rect 57383 8044 57428 8072
rect 56137 8035 56195 8041
rect 57422 8032 57428 8044
rect 57480 8032 57486 8084
rect 54754 7964 54760 8016
rect 54812 8004 54818 8016
rect 55122 8004 55128 8016
rect 54812 7976 55128 8004
rect 54812 7964 54818 7976
rect 55122 7964 55128 7976
rect 55180 8004 55186 8016
rect 55858 8004 55864 8016
rect 55180 7976 55864 8004
rect 55180 7964 55186 7976
rect 55858 7964 55864 7976
rect 55916 7964 55922 8016
rect 55953 8007 56011 8013
rect 55953 7973 55965 8007
rect 55999 8004 56011 8007
rect 55999 7976 56180 8004
rect 55999 7973 56011 7976
rect 55953 7967 56011 7973
rect 54772 7936 54800 7964
rect 56152 7948 56180 7976
rect 54680 7908 54800 7936
rect 54573 7871 54631 7877
rect 54573 7837 54585 7871
rect 54619 7837 54631 7871
rect 54573 7831 54631 7837
rect 54680 7800 54708 7908
rect 54846 7896 54852 7948
rect 54904 7936 54910 7948
rect 56045 7939 56103 7945
rect 56045 7936 56057 7939
rect 54904 7908 56057 7936
rect 54904 7896 54910 7908
rect 56045 7905 56057 7908
rect 56091 7905 56103 7939
rect 56045 7899 56103 7905
rect 56134 7896 56140 7948
rect 56192 7896 56198 7948
rect 54754 7828 54760 7880
rect 54812 7868 54818 7880
rect 55493 7871 55551 7877
rect 55493 7868 55505 7871
rect 54812 7840 55505 7868
rect 54812 7828 54818 7840
rect 55493 7837 55505 7840
rect 55539 7837 55551 7871
rect 55493 7831 55551 7837
rect 55858 7828 55864 7880
rect 55916 7868 55922 7880
rect 56778 7868 56784 7880
rect 55916 7840 56784 7868
rect 55916 7828 55922 7840
rect 56778 7828 56784 7840
rect 56836 7828 56842 7880
rect 53760 7772 54708 7800
rect 49786 7732 49792 7744
rect 47688 7704 49792 7732
rect 46532 7692 46538 7704
rect 49786 7692 49792 7704
rect 49844 7692 49850 7744
rect 51074 7692 51080 7744
rect 51132 7732 51138 7744
rect 51626 7732 51632 7744
rect 51132 7704 51632 7732
rect 51132 7692 51138 7704
rect 51626 7692 51632 7704
rect 51684 7692 51690 7744
rect 52638 7692 52644 7744
rect 52696 7732 52702 7744
rect 54481 7735 54539 7741
rect 54481 7732 54493 7735
rect 52696 7704 54493 7732
rect 52696 7692 52702 7704
rect 54481 7701 54493 7704
rect 54527 7701 54539 7735
rect 54481 7695 54539 7701
rect 55674 7692 55680 7744
rect 55732 7732 55738 7744
rect 56873 7735 56931 7741
rect 56873 7732 56885 7735
rect 55732 7704 56885 7732
rect 55732 7692 55738 7704
rect 56873 7701 56885 7704
rect 56919 7701 56931 7735
rect 57974 7732 57980 7744
rect 57935 7704 57980 7732
rect 56873 7695 56931 7701
rect 57974 7692 57980 7704
rect 58032 7692 58038 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 24765 7531 24823 7537
rect 24765 7497 24777 7531
rect 24811 7528 24823 7531
rect 25777 7531 25835 7537
rect 24811 7500 25728 7528
rect 24811 7497 24823 7500
rect 24765 7491 24823 7497
rect 23842 7420 23848 7472
rect 23900 7460 23906 7472
rect 25406 7460 25412 7472
rect 23900 7432 25412 7460
rect 23900 7420 23906 7432
rect 24688 7401 24716 7432
rect 25406 7420 25412 7432
rect 25464 7420 25470 7472
rect 25700 7460 25728 7500
rect 25777 7497 25789 7531
rect 25823 7528 25835 7531
rect 25866 7528 25872 7540
rect 25823 7500 25872 7528
rect 25823 7497 25835 7500
rect 25777 7491 25835 7497
rect 25866 7488 25872 7500
rect 25924 7488 25930 7540
rect 27062 7488 27068 7540
rect 27120 7528 27126 7540
rect 27157 7531 27215 7537
rect 27157 7528 27169 7531
rect 27120 7500 27169 7528
rect 27120 7488 27126 7500
rect 27157 7497 27169 7500
rect 27203 7497 27215 7531
rect 30285 7531 30343 7537
rect 27157 7491 27215 7497
rect 27448 7500 28120 7528
rect 26970 7460 26976 7472
rect 25700 7432 26976 7460
rect 26970 7420 26976 7432
rect 27028 7460 27034 7472
rect 27448 7460 27476 7500
rect 27028 7432 27476 7460
rect 27028 7420 27034 7432
rect 24673 7395 24731 7401
rect 24673 7361 24685 7395
rect 24719 7361 24731 7395
rect 24946 7392 24952 7404
rect 24907 7364 24952 7392
rect 24673 7355 24731 7361
rect 24946 7352 24952 7364
rect 25004 7352 25010 7404
rect 25958 7392 25964 7404
rect 25919 7364 25964 7392
rect 25958 7352 25964 7364
rect 26016 7352 26022 7404
rect 26053 7395 26111 7401
rect 26053 7361 26065 7395
rect 26099 7361 26111 7395
rect 26234 7392 26240 7404
rect 26195 7364 26240 7392
rect 26053 7355 26111 7361
rect 26068 7324 26096 7355
rect 26234 7352 26240 7364
rect 26292 7352 26298 7404
rect 26326 7352 26332 7404
rect 26384 7392 26390 7404
rect 27341 7395 27399 7401
rect 27341 7392 27353 7395
rect 26384 7364 27353 7392
rect 26384 7352 26390 7364
rect 26988 7336 27016 7364
rect 27341 7361 27353 7364
rect 27387 7361 27399 7395
rect 27341 7355 27399 7361
rect 27614 7352 27620 7404
rect 27672 7392 27678 7404
rect 27801 7398 27859 7401
rect 27801 7395 27936 7398
rect 27672 7364 27717 7392
rect 27672 7352 27678 7364
rect 27801 7361 27813 7395
rect 27847 7392 27936 7395
rect 28092 7392 28120 7500
rect 30285 7497 30297 7531
rect 30331 7497 30343 7531
rect 30285 7491 30343 7497
rect 31389 7531 31447 7537
rect 31389 7497 31401 7531
rect 31435 7528 31447 7531
rect 31570 7528 31576 7540
rect 31435 7500 31576 7528
rect 31435 7497 31447 7500
rect 31389 7491 31447 7497
rect 28718 7420 28724 7472
rect 28776 7460 28782 7472
rect 30300 7460 30328 7491
rect 31570 7488 31576 7500
rect 31628 7528 31634 7540
rect 32490 7528 32496 7540
rect 31628 7500 32496 7528
rect 31628 7488 31634 7500
rect 32490 7488 32496 7500
rect 32548 7488 32554 7540
rect 34517 7531 34575 7537
rect 34517 7528 34529 7531
rect 32793 7500 34529 7528
rect 32793 7460 32821 7500
rect 34517 7497 34529 7500
rect 34563 7528 34575 7531
rect 35342 7528 35348 7540
rect 34563 7500 35348 7528
rect 34563 7497 34575 7500
rect 34517 7491 34575 7497
rect 35342 7488 35348 7500
rect 35400 7488 35406 7540
rect 35618 7488 35624 7540
rect 35676 7528 35682 7540
rect 35676 7500 35721 7528
rect 35676 7488 35682 7500
rect 36630 7488 36636 7540
rect 36688 7528 36694 7540
rect 36817 7531 36875 7537
rect 36817 7528 36829 7531
rect 36688 7500 36829 7528
rect 36688 7488 36694 7500
rect 36817 7497 36829 7500
rect 36863 7497 36875 7531
rect 38381 7531 38439 7537
rect 38381 7528 38393 7531
rect 36817 7491 36875 7497
rect 36924 7500 38393 7528
rect 28776 7432 30328 7460
rect 32692 7432 32821 7460
rect 28776 7420 28782 7432
rect 28629 7395 28687 7401
rect 28629 7392 28641 7395
rect 27847 7370 28028 7392
rect 27847 7361 27859 7370
rect 27908 7364 28028 7370
rect 28092 7364 28641 7392
rect 27801 7355 27859 7361
rect 28000 7336 28028 7364
rect 28629 7361 28641 7364
rect 28675 7392 28687 7395
rect 29086 7392 29092 7404
rect 28675 7364 29092 7392
rect 28675 7361 28687 7364
rect 28629 7355 28687 7361
rect 29086 7352 29092 7364
rect 29144 7352 29150 7404
rect 29454 7392 29460 7404
rect 29415 7364 29460 7392
rect 29454 7352 29460 7364
rect 29512 7352 29518 7404
rect 29638 7392 29644 7404
rect 29599 7364 29644 7392
rect 29638 7352 29644 7364
rect 29696 7352 29702 7404
rect 30466 7392 30472 7404
rect 30427 7364 30472 7392
rect 30466 7352 30472 7364
rect 30524 7352 30530 7404
rect 30653 7395 30711 7401
rect 30653 7361 30665 7395
rect 30699 7392 30711 7395
rect 31294 7392 31300 7404
rect 30699 7364 31300 7392
rect 30699 7361 30711 7364
rect 30653 7355 30711 7361
rect 31294 7352 31300 7364
rect 31352 7352 31358 7404
rect 31478 7352 31484 7404
rect 31536 7392 31542 7404
rect 31573 7395 31631 7401
rect 31573 7392 31585 7395
rect 31536 7364 31585 7392
rect 31536 7352 31542 7364
rect 31573 7361 31585 7364
rect 31619 7361 31631 7395
rect 31573 7355 31631 7361
rect 32030 7352 32036 7404
rect 32088 7392 32094 7404
rect 32692 7392 32720 7432
rect 32858 7420 32864 7472
rect 32916 7460 32922 7472
rect 33045 7463 33103 7469
rect 33045 7460 33057 7463
rect 32916 7432 33057 7460
rect 32916 7420 32922 7432
rect 33045 7429 33057 7432
rect 33091 7460 33103 7463
rect 35710 7460 35716 7472
rect 33091 7432 35716 7460
rect 33091 7429 33103 7432
rect 33045 7423 33103 7429
rect 35710 7420 35716 7432
rect 35768 7460 35774 7472
rect 36924 7460 36952 7500
rect 38381 7497 38393 7500
rect 38427 7528 38439 7531
rect 38930 7528 38936 7540
rect 38427 7500 38936 7528
rect 38427 7497 38439 7500
rect 38381 7491 38439 7497
rect 38930 7488 38936 7500
rect 38988 7488 38994 7540
rect 40402 7488 40408 7540
rect 40460 7528 40466 7540
rect 40773 7531 40831 7537
rect 40773 7528 40785 7531
rect 40460 7500 40785 7528
rect 40460 7488 40466 7500
rect 40773 7497 40785 7500
rect 40819 7497 40831 7531
rect 40773 7491 40831 7497
rect 42794 7488 42800 7540
rect 42852 7528 42858 7540
rect 43346 7528 43352 7540
rect 42852 7500 43352 7528
rect 42852 7488 42858 7500
rect 43346 7488 43352 7500
rect 43404 7528 43410 7540
rect 44193 7531 44251 7537
rect 44193 7528 44205 7531
rect 43404 7500 44205 7528
rect 43404 7488 43410 7500
rect 44193 7497 44205 7500
rect 44239 7497 44251 7531
rect 44193 7491 44251 7497
rect 44450 7488 44456 7540
rect 44508 7528 44514 7540
rect 44821 7531 44879 7537
rect 44821 7528 44833 7531
rect 44508 7500 44833 7528
rect 44508 7488 44514 7500
rect 44821 7497 44833 7500
rect 44867 7497 44879 7531
rect 44821 7491 44879 7497
rect 45738 7488 45744 7540
rect 45796 7528 45802 7540
rect 46017 7531 46075 7537
rect 46017 7528 46029 7531
rect 45796 7500 46029 7528
rect 45796 7488 45802 7500
rect 46017 7497 46029 7500
rect 46063 7497 46075 7531
rect 46017 7491 46075 7497
rect 46124 7500 48084 7528
rect 37458 7460 37464 7472
rect 35768 7432 36952 7460
rect 37419 7432 37464 7460
rect 35768 7420 35774 7432
rect 37458 7420 37464 7432
rect 37516 7420 37522 7472
rect 38010 7420 38016 7472
rect 38068 7460 38074 7472
rect 39485 7463 39543 7469
rect 39485 7460 39497 7463
rect 38068 7432 39497 7460
rect 38068 7420 38074 7432
rect 39485 7429 39497 7432
rect 39531 7460 39543 7463
rect 39574 7460 39580 7472
rect 39531 7432 39580 7460
rect 39531 7429 39543 7432
rect 39485 7423 39543 7429
rect 39574 7420 39580 7432
rect 39632 7420 39638 7472
rect 40678 7460 40684 7472
rect 39684 7432 40684 7460
rect 32088 7364 32720 7392
rect 32088 7352 32094 7364
rect 32692 7336 32720 7364
rect 33594 7352 33600 7404
rect 33652 7392 33658 7404
rect 33689 7395 33747 7401
rect 33689 7392 33701 7395
rect 33652 7364 33701 7392
rect 33652 7352 33658 7364
rect 33689 7361 33701 7364
rect 33735 7361 33747 7395
rect 33689 7355 33747 7361
rect 33778 7352 33784 7404
rect 33836 7392 33842 7404
rect 33836 7364 33881 7392
rect 33836 7352 33842 7364
rect 33962 7352 33968 7404
rect 34020 7392 34026 7404
rect 34020 7364 35848 7392
rect 34020 7352 34026 7364
rect 26694 7324 26700 7336
rect 26068 7296 26700 7324
rect 26694 7284 26700 7296
rect 26752 7284 26758 7336
rect 26970 7284 26976 7336
rect 27028 7284 27034 7336
rect 27525 7327 27583 7333
rect 27525 7293 27537 7327
rect 27571 7324 27583 7327
rect 27890 7324 27896 7336
rect 27571 7296 27896 7324
rect 27571 7293 27583 7296
rect 27525 7287 27583 7293
rect 27890 7284 27896 7296
rect 27948 7284 27954 7336
rect 27982 7284 27988 7336
rect 28040 7284 28046 7336
rect 28353 7327 28411 7333
rect 28353 7293 28365 7327
rect 28399 7324 28411 7327
rect 28442 7324 28448 7336
rect 28399 7296 28448 7324
rect 28399 7293 28411 7296
rect 28353 7287 28411 7293
rect 28442 7284 28448 7296
rect 28500 7284 28506 7336
rect 28902 7284 28908 7336
rect 28960 7324 28966 7336
rect 28997 7327 29055 7333
rect 28997 7324 29009 7327
rect 28960 7296 29009 7324
rect 28960 7284 28966 7296
rect 28997 7293 29009 7296
rect 29043 7293 29055 7327
rect 28997 7287 29055 7293
rect 30282 7284 30288 7336
rect 30340 7324 30346 7336
rect 30561 7327 30619 7333
rect 30561 7324 30573 7327
rect 30340 7296 30573 7324
rect 30340 7284 30346 7296
rect 30561 7293 30573 7296
rect 30607 7293 30619 7327
rect 30561 7287 30619 7293
rect 30745 7327 30803 7333
rect 30745 7293 30757 7327
rect 30791 7293 30803 7327
rect 32490 7324 32496 7336
rect 32451 7296 32496 7324
rect 30745 7287 30803 7293
rect 27430 7256 27436 7268
rect 27391 7228 27436 7256
rect 27430 7216 27436 7228
rect 27488 7216 27494 7268
rect 30098 7256 30104 7268
rect 27632 7228 30104 7256
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 25130 7188 25136 7200
rect 24995 7160 25136 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25130 7148 25136 7160
rect 25188 7148 25194 7200
rect 26234 7148 26240 7200
rect 26292 7188 26298 7200
rect 27632 7188 27660 7228
rect 30098 7216 30104 7228
rect 30156 7216 30162 7268
rect 30190 7216 30196 7268
rect 30248 7256 30254 7268
rect 30760 7256 30788 7287
rect 32490 7284 32496 7296
rect 32548 7284 32554 7336
rect 32674 7324 32680 7336
rect 32587 7296 32680 7324
rect 32674 7284 32680 7296
rect 32732 7284 32738 7336
rect 32766 7284 32772 7336
rect 32824 7324 32830 7336
rect 35161 7327 35219 7333
rect 32824 7296 33824 7324
rect 32824 7284 32830 7296
rect 30248 7228 30788 7256
rect 30248 7216 30254 7228
rect 30834 7216 30840 7268
rect 30892 7256 30898 7268
rect 32907 7259 32965 7265
rect 32907 7256 32919 7259
rect 30892 7228 32919 7256
rect 30892 7216 30898 7228
rect 32907 7225 32919 7228
rect 32953 7256 32965 7259
rect 33686 7256 33692 7268
rect 32953 7228 33692 7256
rect 32953 7225 32965 7228
rect 32907 7219 32965 7225
rect 33686 7216 33692 7228
rect 33744 7216 33750 7268
rect 26292 7160 27660 7188
rect 26292 7148 26298 7160
rect 27706 7148 27712 7200
rect 27764 7188 27770 7200
rect 31662 7188 31668 7200
rect 27764 7160 31668 7188
rect 27764 7148 27770 7160
rect 31662 7148 31668 7160
rect 31720 7148 31726 7200
rect 32769 7191 32827 7197
rect 32769 7157 32781 7191
rect 32815 7188 32827 7191
rect 33226 7188 33232 7200
rect 32815 7160 33232 7188
rect 32815 7157 32827 7160
rect 32769 7151 32827 7157
rect 33226 7148 33232 7160
rect 33284 7148 33290 7200
rect 33502 7188 33508 7200
rect 33463 7160 33508 7188
rect 33502 7148 33508 7160
rect 33560 7148 33566 7200
rect 33796 7188 33824 7296
rect 35161 7293 35173 7327
rect 35207 7324 35219 7327
rect 35342 7324 35348 7336
rect 35207 7296 35348 7324
rect 35207 7293 35219 7296
rect 35161 7287 35219 7293
rect 35342 7284 35348 7296
rect 35400 7284 35406 7336
rect 35820 7324 35848 7364
rect 35894 7352 35900 7404
rect 35952 7392 35958 7404
rect 36449 7395 36507 7401
rect 36449 7392 36461 7395
rect 35952 7364 36461 7392
rect 35952 7352 35958 7364
rect 36449 7361 36461 7364
rect 36495 7361 36507 7395
rect 36630 7392 36636 7404
rect 36591 7364 36636 7392
rect 36449 7355 36507 7361
rect 36630 7352 36636 7364
rect 36688 7352 36694 7404
rect 38197 7395 38255 7401
rect 38197 7392 38209 7395
rect 37108 7364 38209 7392
rect 36998 7324 37004 7336
rect 35820 7296 37004 7324
rect 36998 7284 37004 7296
rect 37056 7284 37062 7336
rect 37108 7268 37136 7364
rect 38197 7361 38209 7364
rect 38243 7361 38255 7395
rect 38197 7355 38255 7361
rect 38286 7352 38292 7404
rect 38344 7392 38350 7404
rect 38344 7364 38389 7392
rect 38344 7352 38350 7364
rect 38654 7352 38660 7404
rect 38712 7392 38718 7404
rect 39117 7395 39175 7401
rect 39117 7392 39129 7395
rect 38712 7364 39129 7392
rect 38712 7352 38718 7364
rect 39117 7361 39129 7364
rect 39163 7392 39175 7395
rect 39684 7392 39712 7432
rect 40678 7420 40684 7432
rect 40736 7420 40742 7472
rect 43990 7460 43996 7472
rect 43951 7432 43996 7460
rect 43990 7420 43996 7432
rect 44048 7420 44054 7472
rect 46124 7460 46152 7500
rect 46290 7460 46296 7472
rect 44192 7432 46152 7460
rect 46251 7432 46296 7460
rect 44192 7404 44220 7432
rect 46290 7420 46296 7432
rect 46348 7420 46354 7472
rect 46382 7420 46388 7472
rect 46440 7460 46446 7472
rect 46440 7432 46485 7460
rect 46440 7420 46446 7432
rect 46934 7420 46940 7472
rect 46992 7460 46998 7472
rect 47121 7463 47179 7469
rect 47121 7460 47133 7463
rect 46992 7432 47133 7460
rect 46992 7420 46998 7432
rect 47121 7429 47133 7432
rect 47167 7429 47179 7463
rect 47121 7423 47179 7429
rect 48056 7460 48084 7500
rect 48130 7488 48136 7540
rect 48188 7528 48194 7540
rect 48188 7500 49004 7528
rect 48188 7488 48194 7500
rect 48406 7460 48412 7472
rect 48056 7432 48412 7460
rect 39163 7364 39712 7392
rect 40129 7395 40187 7401
rect 39163 7361 39175 7364
rect 39117 7355 39175 7361
rect 40129 7361 40141 7395
rect 40175 7392 40187 7395
rect 40954 7392 40960 7404
rect 40175 7364 40448 7392
rect 40915 7364 40960 7392
rect 40175 7361 40187 7364
rect 40129 7355 40187 7361
rect 38010 7324 38016 7336
rect 37971 7296 38016 7324
rect 38010 7284 38016 7296
rect 38068 7284 38074 7336
rect 38565 7327 38623 7333
rect 38565 7293 38577 7327
rect 38611 7324 38623 7327
rect 39390 7324 39396 7336
rect 38611 7296 39396 7324
rect 38611 7293 38623 7296
rect 38565 7287 38623 7293
rect 39390 7284 39396 7296
rect 39448 7324 39454 7336
rect 40144 7324 40172 7355
rect 39448 7296 40172 7324
rect 40313 7327 40371 7333
rect 39448 7284 39454 7296
rect 40313 7293 40325 7327
rect 40359 7293 40371 7327
rect 40420 7324 40448 7364
rect 40954 7352 40960 7364
rect 41012 7352 41018 7404
rect 42886 7392 42892 7404
rect 42847 7364 42892 7392
rect 42886 7352 42892 7364
rect 42944 7352 42950 7404
rect 42978 7352 42984 7404
rect 43036 7392 43042 7404
rect 43162 7392 43168 7404
rect 43036 7364 43168 7392
rect 43036 7352 43042 7364
rect 43162 7352 43168 7364
rect 43220 7392 43226 7404
rect 44082 7392 44088 7404
rect 43220 7364 44088 7392
rect 43220 7352 43226 7364
rect 44082 7352 44088 7364
rect 44140 7352 44146 7404
rect 44174 7352 44180 7404
rect 44232 7352 44238 7404
rect 44910 7352 44916 7404
rect 44968 7392 44974 7404
rect 45281 7395 45339 7401
rect 45281 7392 45293 7395
rect 44968 7364 45293 7392
rect 44968 7352 44974 7364
rect 45281 7361 45293 7364
rect 45327 7361 45339 7395
rect 46198 7392 46204 7404
rect 46159 7364 46204 7392
rect 45281 7355 45339 7361
rect 46198 7352 46204 7364
rect 46256 7352 46262 7404
rect 46523 7395 46581 7401
rect 46523 7361 46535 7395
rect 46569 7392 46581 7395
rect 47210 7392 47216 7404
rect 46569 7364 47216 7392
rect 46569 7361 46581 7364
rect 46523 7355 46581 7361
rect 47210 7352 47216 7364
rect 47268 7352 47274 7404
rect 47578 7352 47584 7404
rect 47636 7392 47642 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 47636 7364 47961 7392
rect 47636 7352 47642 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 41141 7327 41199 7333
rect 41141 7324 41153 7327
rect 40420 7296 41153 7324
rect 40313 7287 40371 7293
rect 41141 7293 41153 7296
rect 41187 7293 41199 7327
rect 41141 7287 41199 7293
rect 33873 7259 33931 7265
rect 33873 7225 33885 7259
rect 33919 7256 33931 7259
rect 34146 7256 34152 7268
rect 33919 7228 34152 7256
rect 33919 7225 33931 7228
rect 33873 7219 33931 7225
rect 34146 7216 34152 7228
rect 34204 7216 34210 7268
rect 35526 7216 35532 7268
rect 35584 7256 35590 7268
rect 37090 7256 37096 7268
rect 35584 7228 37096 7256
rect 35584 7216 35590 7228
rect 37090 7216 37096 7228
rect 37148 7216 37154 7268
rect 39945 7259 40003 7265
rect 39945 7256 39957 7259
rect 37200 7228 39957 7256
rect 37200 7188 37228 7228
rect 39945 7225 39957 7228
rect 39991 7225 40003 7259
rect 40328 7256 40356 7287
rect 42518 7284 42524 7336
rect 42576 7324 42582 7336
rect 42797 7327 42855 7333
rect 42797 7324 42809 7327
rect 42576 7296 42809 7324
rect 42576 7284 42582 7296
rect 42797 7293 42809 7296
rect 42843 7293 42855 7327
rect 42797 7287 42855 7293
rect 43073 7327 43131 7333
rect 43073 7293 43085 7327
rect 43119 7324 43131 7327
rect 43438 7324 43444 7336
rect 43119 7296 43444 7324
rect 43119 7293 43131 7296
rect 43073 7287 43131 7293
rect 43438 7284 43444 7296
rect 43496 7324 43502 7336
rect 46382 7324 46388 7336
rect 43496 7296 46388 7324
rect 43496 7284 43502 7296
rect 46382 7284 46388 7296
rect 46440 7284 46446 7336
rect 46661 7327 46719 7333
rect 46661 7293 46673 7327
rect 46707 7324 46719 7327
rect 47765 7327 47823 7333
rect 47765 7324 47777 7327
rect 46707 7296 47777 7324
rect 46707 7293 46719 7296
rect 46661 7287 46719 7293
rect 47765 7293 47777 7296
rect 47811 7293 47823 7327
rect 48056 7324 48084 7432
rect 48406 7420 48412 7432
rect 48464 7420 48470 7472
rect 48976 7404 49004 7500
rect 50062 7488 50068 7540
rect 50120 7528 50126 7540
rect 51353 7531 51411 7537
rect 51353 7528 51365 7531
rect 50120 7500 51365 7528
rect 50120 7488 50126 7500
rect 51353 7497 51365 7500
rect 51399 7497 51411 7531
rect 51353 7491 51411 7497
rect 51534 7488 51540 7540
rect 51592 7528 51598 7540
rect 52546 7528 52552 7540
rect 51592 7500 52552 7528
rect 51592 7488 51598 7500
rect 52546 7488 52552 7500
rect 52604 7488 52610 7540
rect 52730 7488 52736 7540
rect 52788 7528 52794 7540
rect 53009 7531 53067 7537
rect 53009 7528 53021 7531
rect 52788 7500 53021 7528
rect 52788 7488 52794 7500
rect 53009 7497 53021 7500
rect 53055 7497 53067 7531
rect 53926 7528 53932 7540
rect 53009 7491 53067 7497
rect 53576 7500 53932 7528
rect 51258 7420 51264 7472
rect 51316 7460 51322 7472
rect 51905 7463 51963 7469
rect 51905 7460 51917 7463
rect 51316 7432 51917 7460
rect 51316 7420 51322 7432
rect 51905 7429 51917 7432
rect 51951 7429 51963 7463
rect 51905 7423 51963 7429
rect 52273 7463 52331 7469
rect 52273 7429 52285 7463
rect 52319 7460 52331 7463
rect 53576 7460 53604 7500
rect 53926 7488 53932 7500
rect 53984 7488 53990 7540
rect 54202 7528 54208 7540
rect 54163 7500 54208 7528
rect 54202 7488 54208 7500
rect 54260 7488 54266 7540
rect 56597 7531 56655 7537
rect 56597 7497 56609 7531
rect 56643 7528 56655 7531
rect 56778 7528 56784 7540
rect 56643 7500 56784 7528
rect 56643 7497 56655 7500
rect 56597 7491 56655 7497
rect 56778 7488 56784 7500
rect 56836 7488 56842 7540
rect 54110 7460 54116 7472
rect 52319 7432 53604 7460
rect 53668 7432 54116 7460
rect 52319 7429 52331 7432
rect 52273 7423 52331 7429
rect 48133 7395 48191 7401
rect 48133 7361 48145 7395
rect 48179 7392 48191 7395
rect 48590 7392 48596 7404
rect 48179 7364 48596 7392
rect 48179 7361 48191 7364
rect 48133 7355 48191 7361
rect 48590 7352 48596 7364
rect 48648 7352 48654 7404
rect 48777 7395 48835 7401
rect 48777 7361 48789 7395
rect 48823 7392 48835 7395
rect 48866 7392 48872 7404
rect 48823 7364 48872 7392
rect 48823 7361 48835 7364
rect 48777 7355 48835 7361
rect 48866 7352 48872 7364
rect 48924 7352 48930 7404
rect 48958 7352 48964 7404
rect 49016 7392 49022 7404
rect 49697 7395 49755 7401
rect 49697 7392 49709 7395
rect 49016 7364 49709 7392
rect 49016 7352 49022 7364
rect 49697 7361 49709 7364
rect 49743 7361 49755 7395
rect 49697 7355 49755 7361
rect 49786 7352 49792 7404
rect 49844 7392 49850 7404
rect 50985 7395 51043 7401
rect 49844 7364 49889 7392
rect 49844 7352 49850 7364
rect 50985 7361 50997 7395
rect 51031 7392 51043 7395
rect 51350 7392 51356 7404
rect 51031 7364 51356 7392
rect 51031 7361 51043 7364
rect 50985 7355 51043 7361
rect 51350 7352 51356 7364
rect 51408 7352 51414 7404
rect 51445 7395 51503 7401
rect 51445 7361 51457 7395
rect 51491 7392 51503 7395
rect 52178 7392 52184 7404
rect 51491 7364 52184 7392
rect 51491 7361 51503 7364
rect 51445 7355 51503 7361
rect 52178 7352 52184 7364
rect 52236 7352 52242 7404
rect 48225 7327 48283 7333
rect 48225 7324 48237 7327
rect 48056 7296 48237 7324
rect 47765 7287 47823 7293
rect 48225 7293 48237 7296
rect 48271 7293 48283 7327
rect 49602 7324 49608 7336
rect 48225 7287 48283 7293
rect 48792 7296 49464 7324
rect 49563 7296 49608 7324
rect 40494 7256 40500 7268
rect 40328 7228 40500 7256
rect 39945 7219 40003 7225
rect 33796 7160 37228 7188
rect 37458 7148 37464 7200
rect 37516 7188 37522 7200
rect 38562 7188 38568 7200
rect 37516 7160 38568 7188
rect 37516 7148 37522 7160
rect 38562 7148 38568 7160
rect 38620 7148 38626 7200
rect 39960 7188 39988 7219
rect 40494 7216 40500 7228
rect 40552 7216 40558 7268
rect 40678 7216 40684 7268
rect 40736 7256 40742 7268
rect 41601 7259 41659 7265
rect 41601 7256 41613 7259
rect 40736 7228 41613 7256
rect 40736 7216 40742 7228
rect 41601 7225 41613 7228
rect 41647 7225 41659 7259
rect 44266 7256 44272 7268
rect 44179 7228 44272 7256
rect 41601 7219 41659 7225
rect 41046 7188 41052 7200
rect 39960 7160 41052 7188
rect 41046 7148 41052 7160
rect 41104 7148 41110 7200
rect 41966 7148 41972 7200
rect 42024 7188 42030 7200
rect 44192 7197 44220 7228
rect 44266 7216 44272 7228
rect 44324 7256 44330 7268
rect 47854 7256 47860 7268
rect 44324 7228 47860 7256
rect 44324 7216 44330 7228
rect 47854 7216 47860 7228
rect 47912 7256 47918 7268
rect 48792 7256 48820 7296
rect 47912 7228 48820 7256
rect 48869 7259 48927 7265
rect 47912 7216 47918 7228
rect 48869 7225 48881 7259
rect 48915 7256 48927 7259
rect 49326 7256 49332 7268
rect 48915 7228 49332 7256
rect 48915 7225 48927 7228
rect 48869 7219 48927 7225
rect 49326 7216 49332 7228
rect 49384 7216 49390 7268
rect 49436 7256 49464 7296
rect 49602 7284 49608 7296
rect 49660 7284 49666 7336
rect 49878 7324 49884 7336
rect 49839 7296 49884 7324
rect 49878 7284 49884 7296
rect 49936 7284 49942 7336
rect 51074 7284 51080 7336
rect 51132 7324 51138 7336
rect 52288 7324 52316 7423
rect 52914 7392 52920 7404
rect 52875 7364 52920 7392
rect 52914 7352 52920 7364
rect 52972 7352 52978 7404
rect 53193 7395 53251 7401
rect 53193 7361 53205 7395
rect 53239 7392 53251 7395
rect 53466 7392 53472 7404
rect 53239 7364 53472 7392
rect 53239 7361 53251 7364
rect 53193 7355 53251 7361
rect 53466 7352 53472 7364
rect 53524 7392 53530 7404
rect 53668 7392 53696 7432
rect 54110 7420 54116 7432
rect 54168 7460 54174 7472
rect 56134 7460 56140 7472
rect 54168 7432 56140 7460
rect 54168 7420 54174 7432
rect 54680 7404 54708 7432
rect 56134 7420 56140 7432
rect 56192 7420 56198 7472
rect 53524 7364 53696 7392
rect 53524 7352 53530 7364
rect 53926 7352 53932 7404
rect 53984 7392 53990 7404
rect 54478 7392 54484 7404
rect 53984 7364 54484 7392
rect 53984 7352 53990 7364
rect 54478 7352 54484 7364
rect 54536 7352 54542 7404
rect 54662 7352 54668 7404
rect 54720 7392 54726 7404
rect 54720 7364 54813 7392
rect 54720 7352 54726 7364
rect 54846 7352 54852 7404
rect 54904 7392 54910 7404
rect 58066 7392 58072 7404
rect 54904 7364 54949 7392
rect 58027 7364 58072 7392
rect 54904 7352 54910 7364
rect 58066 7352 58072 7364
rect 58124 7352 58130 7404
rect 51132 7296 51177 7324
rect 51276 7296 52316 7324
rect 51132 7284 51138 7296
rect 51169 7259 51227 7265
rect 49436 7228 51120 7256
rect 42613 7191 42671 7197
rect 42613 7188 42625 7191
rect 42024 7160 42625 7188
rect 42024 7148 42030 7160
rect 42613 7157 42625 7160
rect 42659 7157 42671 7191
rect 42613 7151 42671 7157
rect 44177 7191 44235 7197
rect 44177 7157 44189 7191
rect 44223 7157 44235 7191
rect 44358 7188 44364 7200
rect 44319 7160 44364 7188
rect 44177 7151 44235 7157
rect 44358 7148 44364 7160
rect 44416 7148 44422 7200
rect 45189 7191 45247 7197
rect 45189 7157 45201 7191
rect 45235 7188 45247 7191
rect 45278 7188 45284 7200
rect 45235 7160 45284 7188
rect 45235 7157 45247 7160
rect 45189 7151 45247 7157
rect 45278 7148 45284 7160
rect 45336 7188 45342 7200
rect 47026 7188 47032 7200
rect 45336 7160 47032 7188
rect 45336 7148 45342 7160
rect 47026 7148 47032 7160
rect 47084 7148 47090 7200
rect 49418 7188 49424 7200
rect 49379 7160 49424 7188
rect 49418 7148 49424 7160
rect 49476 7148 49482 7200
rect 49786 7148 49792 7200
rect 49844 7188 49850 7200
rect 50709 7191 50767 7197
rect 50709 7188 50721 7191
rect 49844 7160 50721 7188
rect 49844 7148 49850 7160
rect 50709 7157 50721 7160
rect 50755 7157 50767 7191
rect 51092 7188 51120 7228
rect 51169 7225 51181 7259
rect 51215 7256 51227 7259
rect 51276 7256 51304 7296
rect 53282 7284 53288 7336
rect 53340 7324 53346 7336
rect 54294 7324 54300 7336
rect 53340 7296 54300 7324
rect 53340 7284 53346 7296
rect 54294 7284 54300 7296
rect 54352 7324 54358 7336
rect 54573 7327 54631 7333
rect 54573 7324 54585 7327
rect 54352 7296 54585 7324
rect 54352 7284 54358 7296
rect 54573 7293 54585 7296
rect 54619 7293 54631 7327
rect 54573 7287 54631 7293
rect 56962 7256 56968 7268
rect 51215 7228 51304 7256
rect 51368 7228 56968 7256
rect 51215 7225 51227 7228
rect 51169 7219 51227 7225
rect 51368 7188 51396 7228
rect 56962 7216 56968 7228
rect 57020 7216 57026 7268
rect 51092 7160 51396 7188
rect 50709 7151 50767 7157
rect 51718 7148 51724 7200
rect 51776 7188 51782 7200
rect 52730 7188 52736 7200
rect 51776 7160 52736 7188
rect 51776 7148 51782 7160
rect 52730 7148 52736 7160
rect 52788 7148 52794 7200
rect 53374 7188 53380 7200
rect 53335 7160 53380 7188
rect 53374 7148 53380 7160
rect 53432 7148 53438 7200
rect 53650 7148 53656 7200
rect 53708 7188 53714 7200
rect 54754 7188 54760 7200
rect 53708 7160 54760 7188
rect 53708 7148 53714 7160
rect 54754 7148 54760 7160
rect 54812 7148 54818 7200
rect 55490 7188 55496 7200
rect 55451 7160 55496 7188
rect 55490 7148 55496 7160
rect 55548 7188 55554 7200
rect 55674 7188 55680 7200
rect 55548 7160 55680 7188
rect 55548 7148 55554 7160
rect 55674 7148 55680 7160
rect 55732 7188 55738 7200
rect 55953 7191 56011 7197
rect 55953 7188 55965 7191
rect 55732 7160 55965 7188
rect 55732 7148 55738 7160
rect 55953 7157 55965 7160
rect 55999 7157 56011 7191
rect 55953 7151 56011 7157
rect 56318 7148 56324 7200
rect 56376 7188 56382 7200
rect 57057 7191 57115 7197
rect 57057 7188 57069 7191
rect 56376 7160 57069 7188
rect 56376 7148 56382 7160
rect 57057 7157 57069 7160
rect 57103 7157 57115 7191
rect 57057 7151 57115 7157
rect 57882 7148 57888 7200
rect 57940 7188 57946 7200
rect 58253 7191 58311 7197
rect 58253 7188 58265 7191
rect 57940 7160 58265 7188
rect 57940 7148 57946 7160
rect 58253 7157 58265 7160
rect 58299 7157 58311 7191
rect 58253 7151 58311 7157
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 26789 6987 26847 6993
rect 26789 6953 26801 6987
rect 26835 6984 26847 6987
rect 27430 6984 27436 6996
rect 26835 6956 27436 6984
rect 26835 6953 26847 6956
rect 26789 6947 26847 6953
rect 27430 6944 27436 6956
rect 27488 6944 27494 6996
rect 27614 6944 27620 6996
rect 27672 6984 27678 6996
rect 28077 6987 28135 6993
rect 28077 6984 28089 6987
rect 27672 6956 28089 6984
rect 27672 6944 27678 6956
rect 28077 6953 28089 6956
rect 28123 6953 28135 6987
rect 28077 6947 28135 6953
rect 28350 6944 28356 6996
rect 28408 6984 28414 6996
rect 30834 6984 30840 6996
rect 28408 6956 30840 6984
rect 28408 6944 28414 6956
rect 30834 6944 30840 6956
rect 30892 6944 30898 6996
rect 33781 6987 33839 6993
rect 33781 6953 33793 6987
rect 33827 6984 33839 6987
rect 34054 6984 34060 6996
rect 33827 6956 34060 6984
rect 33827 6953 33839 6956
rect 33781 6947 33839 6953
rect 34054 6944 34060 6956
rect 34112 6944 34118 6996
rect 34146 6944 34152 6996
rect 34204 6984 34210 6996
rect 34790 6984 34796 6996
rect 34204 6956 34796 6984
rect 34204 6944 34210 6956
rect 34790 6944 34796 6956
rect 34848 6984 34854 6996
rect 34977 6987 35035 6993
rect 34977 6984 34989 6987
rect 34848 6956 34989 6984
rect 34848 6944 34854 6956
rect 34977 6953 34989 6956
rect 35023 6953 35035 6987
rect 34977 6947 35035 6953
rect 35434 6944 35440 6996
rect 35492 6984 35498 6996
rect 38654 6984 38660 6996
rect 35492 6956 38660 6984
rect 35492 6944 35498 6956
rect 38654 6944 38660 6956
rect 38712 6944 38718 6996
rect 41138 6944 41144 6996
rect 41196 6984 41202 6996
rect 41877 6987 41935 6993
rect 41877 6984 41889 6987
rect 41196 6956 41889 6984
rect 41196 6944 41202 6956
rect 41877 6953 41889 6956
rect 41923 6953 41935 6987
rect 41877 6947 41935 6953
rect 43714 6944 43720 6996
rect 43772 6984 43778 6996
rect 43809 6987 43867 6993
rect 43809 6984 43821 6987
rect 43772 6956 43821 6984
rect 43772 6944 43778 6956
rect 43809 6953 43821 6956
rect 43855 6984 43867 6987
rect 45554 6984 45560 6996
rect 43855 6956 45560 6984
rect 43855 6953 43867 6956
rect 43809 6947 43867 6953
rect 45554 6944 45560 6956
rect 45612 6944 45618 6996
rect 45738 6944 45744 6996
rect 45796 6984 45802 6996
rect 46934 6984 46940 6996
rect 45796 6956 46940 6984
rect 45796 6944 45802 6956
rect 46934 6944 46940 6956
rect 46992 6944 46998 6996
rect 47210 6984 47216 6996
rect 47171 6956 47216 6984
rect 47210 6944 47216 6956
rect 47268 6944 47274 6996
rect 48133 6987 48191 6993
rect 48133 6953 48145 6987
rect 48179 6984 48191 6987
rect 48222 6984 48228 6996
rect 48179 6956 48228 6984
rect 48179 6953 48191 6956
rect 48133 6947 48191 6953
rect 48222 6944 48228 6956
rect 48280 6944 48286 6996
rect 48501 6987 48559 6993
rect 48501 6953 48513 6987
rect 48547 6984 48559 6987
rect 48590 6984 48596 6996
rect 48547 6956 48596 6984
rect 48547 6953 48559 6956
rect 48501 6947 48559 6953
rect 48590 6944 48596 6956
rect 48648 6944 48654 6996
rect 49418 6944 49424 6996
rect 49476 6984 49482 6996
rect 49513 6987 49571 6993
rect 49513 6984 49525 6987
rect 49476 6956 49525 6984
rect 49476 6944 49482 6956
rect 49513 6953 49525 6956
rect 49559 6953 49571 6987
rect 50798 6984 50804 6996
rect 49513 6947 49571 6953
rect 49804 6956 50804 6984
rect 24302 6876 24308 6928
rect 24360 6916 24366 6928
rect 27062 6916 27068 6928
rect 24360 6888 27068 6916
rect 24360 6876 24366 6888
rect 27062 6876 27068 6888
rect 27120 6876 27126 6928
rect 27246 6876 27252 6928
rect 27304 6916 27310 6928
rect 27632 6916 27660 6944
rect 27304 6888 27660 6916
rect 27304 6876 27310 6888
rect 28810 6876 28816 6928
rect 28868 6916 28874 6928
rect 29638 6916 29644 6928
rect 28868 6888 29644 6916
rect 28868 6876 28874 6888
rect 29638 6876 29644 6888
rect 29696 6916 29702 6928
rect 31110 6916 31116 6928
rect 29696 6888 31116 6916
rect 29696 6876 29702 6888
rect 31110 6876 31116 6888
rect 31168 6876 31174 6928
rect 33594 6916 33600 6928
rect 33060 6888 33600 6916
rect 25332 6820 27752 6848
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6780 24087 6783
rect 25038 6780 25044 6792
rect 24075 6752 25044 6780
rect 24075 6749 24087 6752
rect 24029 6743 24087 6749
rect 25038 6740 25044 6752
rect 25096 6740 25102 6792
rect 25130 6740 25136 6792
rect 25188 6780 25194 6792
rect 25332 6789 25360 6820
rect 25317 6783 25375 6789
rect 25188 6752 25233 6780
rect 25188 6740 25194 6752
rect 25317 6749 25329 6783
rect 25363 6749 25375 6783
rect 25317 6743 25375 6749
rect 25547 6783 25605 6789
rect 25547 6749 25559 6783
rect 25593 6780 25605 6783
rect 25866 6780 25872 6792
rect 25593 6752 25872 6780
rect 25593 6749 25605 6752
rect 25547 6743 25605 6749
rect 25866 6740 25872 6752
rect 25924 6740 25930 6792
rect 26326 6780 26332 6792
rect 26068 6752 26332 6780
rect 24946 6672 24952 6724
rect 25004 6712 25010 6724
rect 25409 6715 25467 6721
rect 25409 6712 25421 6715
rect 25004 6684 25421 6712
rect 25004 6672 25010 6684
rect 25409 6681 25421 6684
rect 25455 6712 25467 6715
rect 26068 6712 26096 6752
rect 26326 6740 26332 6752
rect 26384 6740 26390 6792
rect 26513 6783 26571 6789
rect 26513 6749 26525 6783
rect 26559 6780 26571 6783
rect 26694 6780 26700 6792
rect 26559 6752 26700 6780
rect 26559 6749 26571 6752
rect 26513 6743 26571 6749
rect 26694 6740 26700 6752
rect 26752 6740 26758 6792
rect 27341 6783 27399 6789
rect 27341 6780 27353 6783
rect 27172 6752 27353 6780
rect 25455 6684 26096 6712
rect 25455 6681 25467 6684
rect 25409 6675 25467 6681
rect 26142 6672 26148 6724
rect 26200 6712 26206 6724
rect 26605 6715 26663 6721
rect 26605 6712 26617 6715
rect 26200 6684 26617 6712
rect 26200 6672 26206 6684
rect 26605 6681 26617 6684
rect 26651 6681 26663 6715
rect 26786 6712 26792 6724
rect 26747 6684 26792 6712
rect 26605 6675 26663 6681
rect 25498 6604 25504 6656
rect 25556 6644 25562 6656
rect 25685 6647 25743 6653
rect 25685 6644 25697 6647
rect 25556 6616 25697 6644
rect 25556 6604 25562 6616
rect 25685 6613 25697 6616
rect 25731 6613 25743 6647
rect 26620 6644 26648 6675
rect 26786 6672 26792 6684
rect 26844 6672 26850 6724
rect 27172 6644 27200 6752
rect 27341 6749 27353 6752
rect 27387 6780 27399 6783
rect 27430 6780 27436 6792
rect 27387 6752 27436 6780
rect 27387 6749 27399 6752
rect 27341 6743 27399 6749
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 27522 6740 27528 6792
rect 27580 6780 27586 6792
rect 27580 6752 27625 6780
rect 27580 6740 27586 6752
rect 27246 6672 27252 6724
rect 27304 6712 27310 6724
rect 27304 6684 27349 6712
rect 27304 6672 27310 6684
rect 26620 6616 27200 6644
rect 27724 6644 27752 6820
rect 28074 6808 28080 6860
rect 28132 6848 28138 6860
rect 28261 6851 28319 6857
rect 28261 6848 28273 6851
rect 28132 6820 28273 6848
rect 28132 6808 28138 6820
rect 28261 6817 28273 6820
rect 28307 6848 28319 6851
rect 28307 6820 28488 6848
rect 28307 6817 28319 6820
rect 28261 6811 28319 6817
rect 28460 6792 28488 6820
rect 28534 6808 28540 6860
rect 28592 6848 28598 6860
rect 29822 6848 29828 6860
rect 28592 6820 29828 6848
rect 28592 6808 28598 6820
rect 29822 6808 29828 6820
rect 29880 6808 29886 6860
rect 30190 6808 30196 6860
rect 30248 6848 30254 6860
rect 30285 6851 30343 6857
rect 30285 6848 30297 6851
rect 30248 6820 30297 6848
rect 30248 6808 30254 6820
rect 30285 6817 30297 6820
rect 30331 6817 30343 6851
rect 30285 6811 30343 6817
rect 30653 6851 30711 6857
rect 30653 6817 30665 6851
rect 30699 6848 30711 6851
rect 31386 6848 31392 6860
rect 30699 6820 31392 6848
rect 30699 6817 30711 6820
rect 30653 6811 30711 6817
rect 31386 6808 31392 6820
rect 31444 6808 31450 6860
rect 33060 6857 33088 6888
rect 33594 6876 33600 6888
rect 33652 6916 33658 6928
rect 34698 6916 34704 6928
rect 33652 6888 34704 6916
rect 33652 6876 33658 6888
rect 34698 6876 34704 6888
rect 34756 6876 34762 6928
rect 35069 6919 35127 6925
rect 35069 6885 35081 6919
rect 35115 6916 35127 6919
rect 35618 6916 35624 6928
rect 35115 6888 35624 6916
rect 35115 6885 35127 6888
rect 35069 6879 35127 6885
rect 35618 6876 35624 6888
rect 35676 6876 35682 6928
rect 38286 6916 38292 6928
rect 36280 6888 38292 6916
rect 33045 6851 33103 6857
rect 33045 6848 33057 6851
rect 31864 6820 33057 6848
rect 31864 6792 31892 6820
rect 33045 6817 33057 6820
rect 33091 6817 33103 6851
rect 33045 6811 33103 6817
rect 33137 6851 33195 6857
rect 33137 6817 33149 6851
rect 33183 6848 33195 6851
rect 34054 6848 34060 6860
rect 33183 6820 34060 6848
rect 33183 6817 33195 6820
rect 33137 6811 33195 6817
rect 34054 6808 34060 6820
rect 34112 6808 34118 6860
rect 34149 6851 34207 6857
rect 34149 6817 34161 6851
rect 34195 6848 34207 6851
rect 34238 6848 34244 6860
rect 34195 6820 34244 6848
rect 34195 6817 34207 6820
rect 34149 6811 34207 6817
rect 28350 6780 28356 6792
rect 28311 6752 28356 6780
rect 28350 6740 28356 6752
rect 28408 6740 28414 6792
rect 28442 6740 28448 6792
rect 28500 6780 28506 6792
rect 29181 6783 29239 6789
rect 28500 6752 29132 6780
rect 28500 6740 28506 6752
rect 27798 6672 27804 6724
rect 27856 6712 27862 6724
rect 28077 6715 28135 6721
rect 28077 6712 28089 6715
rect 27856 6684 28089 6712
rect 27856 6672 27862 6684
rect 28077 6681 28089 6684
rect 28123 6681 28135 6715
rect 29104 6712 29132 6752
rect 29181 6749 29193 6783
rect 29227 6780 29239 6783
rect 29638 6780 29644 6792
rect 29227 6752 29644 6780
rect 29227 6749 29239 6752
rect 29181 6743 29239 6749
rect 29638 6740 29644 6752
rect 29696 6780 29702 6792
rect 30469 6783 30527 6789
rect 30469 6780 30481 6783
rect 29696 6752 30481 6780
rect 29696 6740 29702 6752
rect 30469 6749 30481 6752
rect 30515 6749 30527 6783
rect 30469 6743 30527 6749
rect 30374 6712 30380 6724
rect 29104 6684 30380 6712
rect 28077 6675 28135 6681
rect 30374 6672 30380 6684
rect 30432 6672 30438 6724
rect 28537 6647 28595 6653
rect 28537 6644 28549 6647
rect 27724 6616 28549 6644
rect 25685 6607 25743 6613
rect 28537 6613 28549 6616
rect 28583 6644 28595 6647
rect 29914 6644 29920 6656
rect 28583 6616 29920 6644
rect 28583 6613 28595 6616
rect 28537 6607 28595 6613
rect 29914 6604 29920 6616
rect 29972 6604 29978 6656
rect 30484 6644 30512 6743
rect 30558 6740 30564 6792
rect 30616 6780 30622 6792
rect 30745 6783 30803 6789
rect 30745 6780 30757 6783
rect 30616 6752 30757 6780
rect 30616 6740 30622 6752
rect 30745 6749 30757 6752
rect 30791 6749 30803 6783
rect 30745 6743 30803 6749
rect 30837 6783 30895 6789
rect 30837 6749 30849 6783
rect 30883 6749 30895 6783
rect 31018 6780 31024 6792
rect 30979 6752 31024 6780
rect 30837 6743 30895 6749
rect 30852 6712 30880 6743
rect 31018 6740 31024 6752
rect 31076 6740 31082 6792
rect 31110 6740 31116 6792
rect 31168 6780 31174 6792
rect 31481 6783 31539 6789
rect 31481 6780 31493 6783
rect 31168 6752 31493 6780
rect 31168 6740 31174 6752
rect 31481 6749 31493 6752
rect 31527 6749 31539 6783
rect 31846 6780 31852 6792
rect 31759 6752 31852 6780
rect 31481 6743 31539 6749
rect 31846 6740 31852 6752
rect 31904 6740 31910 6792
rect 31941 6783 31999 6789
rect 31941 6749 31953 6783
rect 31987 6780 31999 6783
rect 32122 6780 32128 6792
rect 31987 6752 32128 6780
rect 31987 6749 31999 6752
rect 31941 6743 31999 6749
rect 32122 6740 32128 6752
rect 32180 6740 32186 6792
rect 32674 6780 32680 6792
rect 32636 6752 32680 6780
rect 32674 6740 32680 6752
rect 32732 6740 32738 6792
rect 32769 6783 32827 6789
rect 32769 6749 32781 6783
rect 32815 6779 32827 6783
rect 33502 6780 33508 6792
rect 32876 6779 33508 6780
rect 32815 6752 33508 6779
rect 32815 6751 32904 6752
rect 32815 6749 32827 6751
rect 32769 6743 32827 6749
rect 33502 6740 33508 6752
rect 33560 6740 33566 6792
rect 33594 6740 33600 6792
rect 33652 6780 33658 6792
rect 33870 6780 33876 6792
rect 33652 6752 33876 6780
rect 33652 6740 33658 6752
rect 33870 6740 33876 6752
rect 33928 6780 33934 6792
rect 33965 6783 34023 6789
rect 33965 6780 33977 6783
rect 33928 6752 33977 6780
rect 33928 6740 33934 6752
rect 33965 6749 33977 6752
rect 34011 6749 34023 6783
rect 33965 6743 34023 6749
rect 30852 6684 32628 6712
rect 31662 6644 31668 6656
rect 30484 6616 31668 6644
rect 31662 6604 31668 6616
rect 31720 6604 31726 6656
rect 31772 6653 31800 6684
rect 31757 6647 31815 6653
rect 31757 6613 31769 6647
rect 31803 6644 31815 6647
rect 32490 6644 32496 6656
rect 31803 6616 31837 6644
rect 32451 6616 32496 6644
rect 31803 6613 31815 6616
rect 31757 6607 31815 6613
rect 32490 6604 32496 6616
rect 32548 6604 32554 6656
rect 32600 6644 32628 6684
rect 33134 6672 33140 6724
rect 33192 6712 33198 6724
rect 34164 6712 34192 6811
rect 34238 6808 34244 6820
rect 34296 6808 34302 6860
rect 35437 6851 35495 6857
rect 35437 6817 35449 6851
rect 35483 6848 35495 6851
rect 35710 6848 35716 6860
rect 35483 6820 35716 6848
rect 35483 6817 35495 6820
rect 35437 6811 35495 6817
rect 35710 6808 35716 6820
rect 35768 6808 35774 6860
rect 35894 6780 35900 6792
rect 33192 6684 34192 6712
rect 34256 6752 35900 6780
rect 33192 6672 33198 6684
rect 34256 6644 34284 6752
rect 35894 6740 35900 6752
rect 35952 6740 35958 6792
rect 36078 6780 36084 6792
rect 36039 6752 36084 6780
rect 36078 6740 36084 6752
rect 36136 6740 36142 6792
rect 36170 6740 36176 6792
rect 36228 6780 36234 6792
rect 36280 6789 36308 6888
rect 38286 6876 38292 6888
rect 38344 6876 38350 6928
rect 41325 6919 41383 6925
rect 41325 6885 41337 6919
rect 41371 6916 41383 6919
rect 41598 6916 41604 6928
rect 41371 6888 41604 6916
rect 41371 6885 41383 6888
rect 41325 6879 41383 6885
rect 41598 6876 41604 6888
rect 41656 6876 41662 6928
rect 43622 6876 43628 6928
rect 43680 6916 43686 6928
rect 46477 6919 46535 6925
rect 46477 6916 46489 6919
rect 43680 6888 46489 6916
rect 43680 6876 43686 6888
rect 46477 6885 46489 6888
rect 46523 6916 46535 6919
rect 46566 6916 46572 6928
rect 46523 6888 46572 6916
rect 46523 6885 46535 6888
rect 46477 6879 46535 6885
rect 46566 6876 46572 6888
rect 46624 6876 46630 6928
rect 46658 6876 46664 6928
rect 46716 6916 46722 6928
rect 49804 6916 49832 6956
rect 50798 6944 50804 6956
rect 50856 6944 50862 6996
rect 52914 6984 52920 6996
rect 51184 6956 52920 6984
rect 46716 6888 47440 6916
rect 46716 6876 46722 6888
rect 47412 6860 47440 6888
rect 48608 6888 49832 6916
rect 37093 6851 37151 6857
rect 37093 6817 37105 6851
rect 37139 6848 37151 6851
rect 37182 6848 37188 6860
rect 37139 6820 37188 6848
rect 37139 6817 37151 6820
rect 37093 6811 37151 6817
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 41966 6848 41972 6860
rect 41156 6820 41972 6848
rect 36265 6783 36323 6789
rect 36265 6780 36277 6783
rect 36228 6752 36277 6780
rect 36228 6740 36234 6752
rect 36265 6749 36277 6752
rect 36311 6749 36323 6783
rect 36265 6743 36323 6749
rect 37553 6783 37611 6789
rect 37553 6749 37565 6783
rect 37599 6780 37611 6783
rect 37642 6780 37648 6792
rect 37599 6752 37648 6780
rect 37599 6749 37611 6752
rect 37553 6743 37611 6749
rect 37642 6740 37648 6752
rect 37700 6740 37706 6792
rect 38010 6780 38016 6792
rect 37971 6752 38016 6780
rect 38010 6740 38016 6752
rect 38068 6740 38074 6792
rect 39482 6780 39488 6792
rect 39443 6752 39488 6780
rect 39482 6740 39488 6752
rect 39540 6740 39546 6792
rect 40218 6780 40224 6792
rect 40179 6752 40224 6780
rect 40218 6740 40224 6752
rect 40276 6740 40282 6792
rect 40494 6740 40500 6792
rect 40552 6780 40558 6792
rect 41156 6789 41184 6820
rect 41966 6808 41972 6820
rect 42024 6808 42030 6860
rect 42518 6848 42524 6860
rect 42479 6820 42524 6848
rect 42518 6808 42524 6820
rect 42576 6808 42582 6860
rect 42886 6848 42892 6860
rect 42812 6820 42892 6848
rect 41141 6783 41199 6789
rect 40552 6752 41092 6780
rect 40552 6740 40558 6752
rect 36096 6712 36124 6740
rect 36722 6712 36728 6724
rect 36096 6684 36728 6712
rect 36722 6672 36728 6684
rect 36780 6672 36786 6724
rect 37734 6672 37740 6724
rect 37792 6712 37798 6724
rect 40957 6715 41015 6721
rect 40957 6712 40969 6715
rect 37792 6684 40969 6712
rect 37792 6672 37798 6684
rect 40957 6681 40969 6684
rect 41003 6681 41015 6715
rect 41064 6712 41092 6752
rect 41141 6749 41153 6783
rect 41187 6749 41199 6783
rect 41414 6780 41420 6792
rect 41375 6752 41420 6780
rect 41141 6743 41199 6749
rect 41414 6740 41420 6752
rect 41472 6740 41478 6792
rect 42613 6783 42671 6789
rect 42613 6749 42625 6783
rect 42659 6780 42671 6783
rect 42812 6780 42840 6820
rect 42886 6808 42892 6820
rect 42944 6808 42950 6860
rect 42981 6851 43039 6857
rect 42981 6817 42993 6851
rect 43027 6848 43039 6851
rect 45370 6848 45376 6860
rect 43027 6820 45376 6848
rect 43027 6817 43039 6820
rect 42981 6811 43039 6817
rect 45370 6808 45376 6820
rect 45428 6808 45434 6860
rect 46750 6848 46756 6860
rect 45480 6820 46756 6848
rect 45480 6789 45508 6820
rect 46750 6808 46756 6820
rect 46808 6808 46814 6860
rect 47394 6848 47400 6860
rect 47307 6820 47400 6848
rect 47394 6808 47400 6820
rect 47452 6808 47458 6860
rect 44453 6783 44511 6789
rect 44453 6780 44465 6783
rect 42659 6752 42840 6780
rect 42904 6752 44465 6780
rect 42659 6749 42671 6752
rect 42613 6743 42671 6749
rect 42904 6712 42932 6752
rect 44453 6749 44465 6752
rect 44499 6749 44511 6783
rect 44453 6743 44511 6749
rect 45465 6783 45523 6789
rect 45465 6749 45477 6783
rect 45511 6749 45523 6783
rect 45465 6743 45523 6749
rect 45833 6783 45891 6789
rect 45833 6749 45845 6783
rect 45879 6780 45891 6783
rect 45879 6752 45968 6780
rect 45879 6749 45891 6752
rect 45833 6743 45891 6749
rect 41064 6684 42932 6712
rect 40957 6675 41015 6681
rect 42978 6672 42984 6724
rect 43036 6712 43042 6724
rect 43898 6712 43904 6724
rect 43036 6684 43760 6712
rect 43859 6684 43904 6712
rect 43036 6672 43042 6684
rect 32600 6616 34284 6644
rect 36265 6647 36323 6653
rect 36265 6613 36277 6647
rect 36311 6644 36323 6647
rect 39114 6644 39120 6656
rect 36311 6616 39120 6644
rect 36311 6613 36323 6616
rect 36265 6607 36323 6613
rect 39114 6604 39120 6616
rect 39172 6604 39178 6656
rect 39298 6644 39304 6656
rect 39259 6616 39304 6644
rect 39298 6604 39304 6616
rect 39356 6604 39362 6656
rect 40402 6644 40408 6656
rect 40315 6616 40408 6644
rect 40402 6604 40408 6616
rect 40460 6644 40466 6656
rect 41414 6644 41420 6656
rect 40460 6616 41420 6644
rect 40460 6604 40466 6616
rect 41414 6604 41420 6616
rect 41472 6604 41478 6656
rect 43732 6644 43760 6684
rect 43898 6672 43904 6684
rect 43956 6672 43962 6724
rect 44358 6672 44364 6724
rect 44416 6712 44422 6724
rect 45278 6712 45284 6724
rect 44416 6684 45284 6712
rect 44416 6672 44422 6684
rect 45278 6672 45284 6684
rect 45336 6712 45342 6724
rect 45649 6715 45707 6721
rect 45649 6712 45661 6715
rect 45336 6684 45661 6712
rect 45336 6672 45342 6684
rect 45649 6681 45661 6684
rect 45695 6681 45707 6715
rect 45649 6675 45707 6681
rect 45738 6672 45744 6724
rect 45796 6712 45802 6724
rect 45940 6712 45968 6752
rect 47302 6740 47308 6792
rect 47360 6780 47366 6792
rect 47578 6780 47584 6792
rect 47360 6752 47405 6780
rect 47539 6752 47584 6780
rect 47360 6740 47366 6752
rect 47578 6740 47584 6752
rect 47636 6740 47642 6792
rect 47670 6740 47676 6792
rect 47728 6780 47734 6792
rect 47728 6752 47773 6780
rect 47728 6740 47734 6752
rect 48038 6740 48044 6792
rect 48096 6780 48102 6792
rect 48608 6789 48636 6888
rect 50154 6876 50160 6928
rect 50212 6916 50218 6928
rect 50433 6919 50491 6925
rect 50433 6916 50445 6919
rect 50212 6888 50445 6916
rect 50212 6876 50218 6888
rect 50433 6885 50445 6888
rect 50479 6916 50491 6919
rect 51184 6916 51212 6956
rect 50479 6888 51212 6916
rect 50479 6885 50491 6888
rect 50433 6879 50491 6885
rect 51258 6876 51264 6928
rect 51316 6916 51322 6928
rect 51316 6888 51856 6916
rect 51316 6876 51322 6888
rect 49050 6848 49056 6860
rect 49011 6820 49056 6848
rect 49050 6808 49056 6820
rect 49108 6808 49114 6860
rect 49786 6848 49792 6860
rect 49252 6820 49792 6848
rect 49252 6789 49280 6820
rect 49786 6808 49792 6820
rect 49844 6808 49850 6860
rect 51828 6857 51856 6888
rect 51813 6851 51871 6857
rect 51813 6817 51825 6851
rect 51859 6817 51871 6851
rect 51813 6811 51871 6817
rect 51920 6792 51948 6956
rect 52914 6944 52920 6956
rect 52972 6944 52978 6996
rect 56318 6984 56324 6996
rect 54462 6956 56324 6984
rect 52822 6876 52828 6928
rect 52880 6916 52886 6928
rect 54462 6916 54490 6956
rect 56318 6944 56324 6956
rect 56376 6944 56382 6996
rect 58066 6984 58072 6996
rect 58027 6956 58072 6984
rect 58066 6944 58072 6956
rect 58124 6944 58130 6996
rect 54662 6916 54668 6928
rect 52880 6888 54490 6916
rect 54623 6888 54668 6916
rect 52880 6876 52886 6888
rect 54662 6876 54668 6888
rect 54720 6876 54726 6928
rect 52454 6848 52460 6860
rect 52196 6820 52460 6848
rect 48593 6783 48651 6789
rect 48593 6780 48605 6783
rect 48096 6752 48605 6780
rect 48096 6740 48102 6752
rect 48593 6749 48605 6752
rect 48639 6749 48651 6783
rect 48593 6743 48651 6749
rect 49237 6783 49295 6789
rect 49237 6749 49249 6783
rect 49283 6749 49295 6783
rect 49237 6743 49295 6749
rect 49326 6740 49332 6792
rect 49384 6780 49390 6792
rect 49605 6783 49663 6789
rect 49384 6752 49429 6780
rect 49384 6740 49390 6752
rect 49605 6749 49617 6783
rect 49651 6780 49663 6783
rect 49878 6780 49884 6792
rect 49651 6752 49884 6780
rect 49651 6749 49663 6752
rect 49605 6743 49663 6749
rect 49878 6740 49884 6752
rect 49936 6740 49942 6792
rect 50338 6780 50344 6792
rect 50299 6752 50344 6780
rect 50338 6740 50344 6752
rect 50396 6740 50402 6792
rect 50609 6783 50667 6789
rect 50609 6749 50621 6783
rect 50655 6782 50667 6783
rect 50798 6782 50804 6792
rect 50655 6754 50804 6782
rect 50655 6749 50667 6754
rect 50609 6743 50667 6749
rect 50798 6740 50804 6754
rect 50856 6740 50862 6792
rect 51718 6780 51724 6792
rect 51679 6752 51724 6780
rect 51718 6740 51724 6752
rect 51776 6740 51782 6792
rect 51902 6740 51908 6792
rect 51960 6780 51966 6792
rect 51960 6752 52053 6780
rect 51960 6740 51966 6752
rect 48682 6712 48688 6724
rect 45796 6684 45841 6712
rect 45940 6684 48688 6712
rect 45796 6672 45802 6684
rect 48682 6672 48688 6684
rect 48740 6672 48746 6724
rect 52196 6712 52224 6820
rect 52454 6808 52460 6820
rect 52512 6808 52518 6860
rect 55214 6808 55220 6860
rect 55272 6848 55278 6860
rect 55493 6851 55551 6857
rect 55493 6848 55505 6851
rect 55272 6820 55505 6848
rect 55272 6808 55278 6820
rect 55493 6817 55505 6820
rect 55539 6817 55551 6851
rect 55493 6811 55551 6817
rect 56226 6808 56232 6860
rect 56284 6848 56290 6860
rect 56873 6851 56931 6857
rect 56873 6848 56885 6851
rect 56284 6820 56885 6848
rect 56284 6808 56290 6820
rect 56873 6817 56885 6820
rect 56919 6817 56931 6851
rect 56873 6811 56931 6817
rect 57330 6808 57336 6860
rect 57388 6848 57394 6860
rect 57425 6851 57483 6857
rect 57425 6848 57437 6851
rect 57388 6820 57437 6848
rect 57388 6808 57394 6820
rect 57425 6817 57437 6820
rect 57471 6817 57483 6851
rect 57425 6811 57483 6817
rect 52270 6740 52276 6792
rect 52328 6780 52334 6792
rect 52549 6783 52607 6789
rect 52549 6780 52561 6783
rect 52328 6752 52561 6780
rect 52328 6740 52334 6752
rect 52549 6749 52561 6752
rect 52595 6749 52607 6783
rect 52549 6743 52607 6749
rect 54754 6740 54760 6792
rect 54812 6780 54818 6792
rect 55677 6783 55735 6789
rect 55677 6780 55689 6783
rect 54812 6752 55689 6780
rect 54812 6740 54818 6752
rect 55677 6749 55689 6752
rect 55723 6749 55735 6783
rect 55677 6743 55735 6749
rect 55769 6783 55827 6789
rect 55769 6749 55781 6783
rect 55815 6749 55827 6783
rect 55769 6743 55827 6749
rect 58253 6783 58311 6789
rect 58253 6749 58265 6783
rect 58299 6780 58311 6783
rect 58526 6780 58532 6792
rect 58299 6752 58532 6780
rect 58299 6749 58311 6752
rect 58253 6743 58311 6749
rect 50816 6684 52224 6712
rect 52365 6715 52423 6721
rect 45922 6644 45928 6656
rect 43732 6616 45928 6644
rect 45922 6604 45928 6616
rect 45980 6604 45986 6656
rect 46017 6647 46075 6653
rect 46017 6613 46029 6647
rect 46063 6644 46075 6647
rect 46290 6644 46296 6656
rect 46063 6616 46296 6644
rect 46063 6613 46075 6616
rect 46017 6607 46075 6613
rect 46290 6604 46296 6616
rect 46348 6604 46354 6656
rect 47394 6604 47400 6656
rect 47452 6644 47458 6656
rect 50816 6653 50844 6684
rect 52365 6681 52377 6715
rect 52411 6712 52423 6715
rect 52454 6712 52460 6724
rect 52411 6684 52460 6712
rect 52411 6681 52423 6684
rect 52365 6675 52423 6681
rect 52454 6672 52460 6684
rect 52512 6672 52518 6724
rect 53282 6712 53288 6724
rect 52564 6684 52868 6712
rect 53243 6684 53288 6712
rect 52564 6656 52592 6684
rect 50801 6647 50859 6653
rect 50801 6644 50813 6647
rect 47452 6616 50813 6644
rect 47452 6604 47458 6616
rect 50801 6613 50813 6616
rect 50847 6613 50859 6647
rect 50801 6607 50859 6613
rect 52546 6604 52552 6656
rect 52604 6604 52610 6656
rect 52730 6644 52736 6656
rect 52691 6616 52736 6644
rect 52730 6604 52736 6616
rect 52788 6604 52794 6656
rect 52840 6644 52868 6684
rect 53282 6672 53288 6684
rect 53340 6672 53346 6724
rect 54846 6712 54852 6724
rect 54807 6684 54852 6712
rect 54846 6672 54852 6684
rect 54904 6712 54910 6724
rect 55030 6712 55036 6724
rect 54904 6684 55036 6712
rect 54904 6672 54910 6684
rect 55030 6672 55036 6684
rect 55088 6672 55094 6724
rect 55784 6712 55812 6743
rect 58526 6740 58532 6752
rect 58584 6740 58590 6792
rect 55692 6684 55812 6712
rect 53377 6647 53435 6653
rect 53377 6644 53389 6647
rect 52840 6616 53389 6644
rect 53377 6613 53389 6616
rect 53423 6644 53435 6647
rect 54110 6644 54116 6656
rect 53423 6616 54116 6644
rect 53423 6613 53435 6616
rect 53377 6607 53435 6613
rect 54110 6604 54116 6616
rect 54168 6604 54174 6656
rect 54202 6604 54208 6656
rect 54260 6644 54266 6656
rect 55692 6644 55720 6684
rect 54260 6616 55720 6644
rect 54260 6604 54266 6616
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 24118 6440 24124 6452
rect 24079 6412 24124 6440
rect 24118 6400 24124 6412
rect 24176 6400 24182 6452
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 27157 6443 27215 6449
rect 27157 6440 27169 6443
rect 25280 6412 27169 6440
rect 25280 6400 25286 6412
rect 27157 6409 27169 6412
rect 27203 6409 27215 6443
rect 28994 6440 29000 6452
rect 28955 6412 29000 6440
rect 27157 6403 27215 6409
rect 28994 6400 29000 6412
rect 29052 6400 29058 6452
rect 29638 6440 29644 6452
rect 29599 6412 29644 6440
rect 29638 6400 29644 6412
rect 29696 6400 29702 6452
rect 29932 6412 30880 6440
rect 24136 6304 24164 6400
rect 25406 6332 25412 6384
rect 25464 6372 25470 6384
rect 25593 6375 25651 6381
rect 25593 6372 25605 6375
rect 25464 6344 25605 6372
rect 25464 6332 25470 6344
rect 25593 6341 25605 6344
rect 25639 6341 25651 6375
rect 25593 6335 25651 6341
rect 28074 6332 28080 6384
rect 28132 6372 28138 6384
rect 28350 6372 28356 6384
rect 28132 6344 28356 6372
rect 28132 6332 28138 6344
rect 28350 6332 28356 6344
rect 28408 6372 28414 6384
rect 29822 6372 29828 6384
rect 28408 6344 29828 6372
rect 28408 6332 28414 6344
rect 24581 6307 24639 6313
rect 24581 6304 24593 6307
rect 24136 6276 24593 6304
rect 24581 6273 24593 6276
rect 24627 6273 24639 6307
rect 25314 6304 25320 6316
rect 25275 6276 25320 6304
rect 24581 6267 24639 6273
rect 25314 6264 25320 6276
rect 25372 6264 25378 6316
rect 25869 6307 25927 6313
rect 25869 6273 25881 6307
rect 25915 6273 25927 6307
rect 26050 6304 26056 6316
rect 26011 6276 26056 6304
rect 25869 6267 25927 6273
rect 24857 6239 24915 6245
rect 24857 6205 24869 6239
rect 24903 6236 24915 6239
rect 25774 6236 25780 6248
rect 24903 6208 25780 6236
rect 24903 6205 24915 6208
rect 24857 6199 24915 6205
rect 25774 6196 25780 6208
rect 25832 6196 25838 6248
rect 25884 6236 25912 6267
rect 26050 6264 26056 6276
rect 26108 6264 26114 6316
rect 28736 6313 28764 6344
rect 29822 6332 29828 6344
rect 29880 6372 29886 6384
rect 29932 6372 29960 6412
rect 30285 6375 30343 6381
rect 30285 6372 30297 6375
rect 29880 6344 29960 6372
rect 30024 6344 30297 6372
rect 29880 6332 29886 6344
rect 28721 6307 28779 6313
rect 28721 6273 28733 6307
rect 28767 6273 28779 6307
rect 28721 6267 28779 6273
rect 26326 6236 26332 6248
rect 25884 6208 26332 6236
rect 26326 6196 26332 6208
rect 26384 6196 26390 6248
rect 26605 6239 26663 6245
rect 26605 6205 26617 6239
rect 26651 6236 26663 6239
rect 26694 6236 26700 6248
rect 26651 6208 26700 6236
rect 26651 6205 26663 6208
rect 26605 6199 26663 6205
rect 26694 6196 26700 6208
rect 26752 6196 26758 6248
rect 27430 6196 27436 6248
rect 27488 6236 27494 6248
rect 28350 6236 28356 6248
rect 27488 6208 28356 6236
rect 27488 6196 27494 6208
rect 28350 6196 28356 6208
rect 28408 6236 28414 6248
rect 30024 6236 30052 6344
rect 30285 6341 30297 6344
rect 30331 6341 30343 6375
rect 30285 6335 30343 6341
rect 30469 6375 30527 6381
rect 30469 6341 30481 6375
rect 30515 6372 30527 6375
rect 30742 6372 30748 6384
rect 30515 6344 30748 6372
rect 30515 6341 30527 6344
rect 30469 6335 30527 6341
rect 30101 6307 30159 6313
rect 30101 6273 30113 6307
rect 30147 6273 30159 6307
rect 30300 6304 30328 6335
rect 30742 6332 30748 6344
rect 30800 6332 30806 6384
rect 30852 6372 30880 6412
rect 30926 6400 30932 6452
rect 30984 6440 30990 6452
rect 31021 6443 31079 6449
rect 31021 6440 31033 6443
rect 30984 6412 31033 6440
rect 30984 6400 30990 6412
rect 31021 6409 31033 6412
rect 31067 6409 31079 6443
rect 31021 6403 31079 6409
rect 31757 6443 31815 6449
rect 31757 6409 31769 6443
rect 31803 6440 31815 6443
rect 32122 6440 32128 6452
rect 31803 6412 32128 6440
rect 31803 6409 31815 6412
rect 31757 6403 31815 6409
rect 32122 6400 32128 6412
rect 32180 6400 32186 6452
rect 32493 6443 32551 6449
rect 32493 6409 32505 6443
rect 32539 6409 32551 6443
rect 32493 6403 32551 6409
rect 31478 6372 31484 6384
rect 30852 6344 31484 6372
rect 30558 6304 30564 6316
rect 30300 6276 30564 6304
rect 30101 6267 30159 6273
rect 28408 6208 30052 6236
rect 30116 6236 30144 6267
rect 30558 6264 30564 6276
rect 30616 6264 30622 6316
rect 30944 6313 30972 6344
rect 31478 6332 31484 6344
rect 31536 6332 31542 6384
rect 32508 6372 32536 6403
rect 32582 6400 32588 6452
rect 32640 6440 32646 6452
rect 33873 6443 33931 6449
rect 33873 6440 33885 6443
rect 32640 6412 33885 6440
rect 32640 6400 32646 6412
rect 33873 6409 33885 6412
rect 33919 6409 33931 6443
rect 33873 6403 33931 6409
rect 34054 6400 34060 6452
rect 34112 6440 34118 6452
rect 39850 6440 39856 6452
rect 34112 6412 39856 6440
rect 34112 6400 34118 6412
rect 39850 6400 39856 6412
rect 39908 6400 39914 6452
rect 40497 6443 40555 6449
rect 40497 6409 40509 6443
rect 40543 6440 40555 6443
rect 40954 6440 40960 6452
rect 40543 6412 40960 6440
rect 40543 6409 40555 6412
rect 40497 6403 40555 6409
rect 32674 6372 32680 6384
rect 32508 6344 32680 6372
rect 32674 6332 32680 6344
rect 32732 6372 32738 6384
rect 33134 6372 33140 6384
rect 32732 6344 33140 6372
rect 32732 6332 32738 6344
rect 33134 6332 33140 6344
rect 33192 6332 33198 6384
rect 33229 6375 33287 6381
rect 33229 6341 33241 6375
rect 33275 6372 33287 6375
rect 33502 6372 33508 6384
rect 33275 6344 33508 6372
rect 33275 6341 33287 6344
rect 33229 6335 33287 6341
rect 33502 6332 33508 6344
rect 33560 6332 33566 6384
rect 34606 6372 34612 6384
rect 34348 6344 34612 6372
rect 30929 6307 30987 6313
rect 30929 6273 30941 6307
rect 30975 6273 30987 6307
rect 30929 6267 30987 6273
rect 31113 6307 31171 6313
rect 31113 6273 31125 6307
rect 31159 6304 31171 6307
rect 31294 6304 31300 6316
rect 31159 6276 31300 6304
rect 31159 6273 31171 6276
rect 31113 6267 31171 6273
rect 31294 6264 31300 6276
rect 31352 6264 31358 6316
rect 31386 6264 31392 6316
rect 31444 6304 31450 6316
rect 32309 6307 32367 6313
rect 32309 6304 32321 6307
rect 31444 6276 32321 6304
rect 31444 6264 31450 6276
rect 32309 6273 32321 6276
rect 32355 6273 32367 6307
rect 33686 6304 33692 6316
rect 33647 6276 33692 6304
rect 32309 6267 32367 6273
rect 33686 6264 33692 6276
rect 33744 6264 33750 6316
rect 34057 6307 34115 6313
rect 34057 6273 34069 6307
rect 34103 6304 34115 6307
rect 34238 6304 34244 6316
rect 34103 6276 34244 6304
rect 34103 6273 34115 6276
rect 34057 6267 34115 6273
rect 34238 6264 34244 6276
rect 34296 6264 34302 6316
rect 34348 6313 34376 6344
rect 34606 6332 34612 6344
rect 34664 6372 34670 6384
rect 36446 6372 36452 6384
rect 34664 6344 36308 6372
rect 36407 6344 36452 6372
rect 34664 6332 34670 6344
rect 34333 6307 34391 6313
rect 34333 6273 34345 6307
rect 34379 6273 34391 6307
rect 34333 6267 34391 6273
rect 35069 6307 35127 6313
rect 35069 6273 35081 6307
rect 35115 6304 35127 6307
rect 35710 6304 35716 6316
rect 35115 6276 35716 6304
rect 35115 6273 35127 6276
rect 35069 6267 35127 6273
rect 35710 6264 35716 6276
rect 35768 6264 35774 6316
rect 36280 6313 36308 6344
rect 36446 6332 36452 6344
rect 36504 6332 36510 6384
rect 38010 6372 38016 6384
rect 36924 6344 38016 6372
rect 36924 6316 36952 6344
rect 38010 6332 38016 6344
rect 38068 6332 38074 6384
rect 38194 6332 38200 6384
rect 38252 6372 38258 6384
rect 38654 6372 38660 6384
rect 38252 6344 38660 6372
rect 38252 6332 38258 6344
rect 38654 6332 38660 6344
rect 38712 6372 38718 6384
rect 38712 6344 38792 6372
rect 38712 6332 38718 6344
rect 36265 6307 36323 6313
rect 36265 6273 36277 6307
rect 36311 6304 36323 6307
rect 36354 6304 36360 6316
rect 36311 6276 36360 6304
rect 36311 6273 36323 6276
rect 36265 6267 36323 6273
rect 36354 6264 36360 6276
rect 36412 6264 36418 6316
rect 36906 6304 36912 6316
rect 36867 6276 36912 6304
rect 36906 6264 36912 6276
rect 36964 6264 36970 6316
rect 37090 6264 37096 6316
rect 37148 6304 37154 6316
rect 37553 6307 37611 6313
rect 37553 6304 37565 6307
rect 37148 6276 37565 6304
rect 37148 6264 37154 6276
rect 37553 6273 37565 6276
rect 37599 6304 37611 6307
rect 38102 6304 38108 6316
rect 37599 6276 38108 6304
rect 37599 6273 37611 6276
rect 37553 6267 37611 6273
rect 38102 6264 38108 6276
rect 38160 6264 38166 6316
rect 38764 6313 38792 6344
rect 38838 6332 38844 6384
rect 38896 6381 38902 6384
rect 38896 6372 38903 6381
rect 38896 6344 38941 6372
rect 38896 6335 38903 6344
rect 38896 6332 38902 6335
rect 38749 6307 38807 6313
rect 38749 6273 38761 6307
rect 38795 6273 38807 6307
rect 38930 6304 38936 6316
rect 38891 6276 38936 6304
rect 38749 6267 38807 6273
rect 38930 6264 38936 6276
rect 38988 6264 38994 6316
rect 39114 6264 39120 6316
rect 39172 6304 39178 6316
rect 39850 6304 39856 6316
rect 39172 6276 39265 6304
rect 39811 6276 39856 6304
rect 39172 6264 39178 6276
rect 30374 6236 30380 6248
rect 30116 6208 30380 6236
rect 28408 6196 28414 6208
rect 30374 6196 30380 6208
rect 30432 6236 30438 6248
rect 33134 6236 33140 6248
rect 30432 6208 33140 6236
rect 30432 6196 30438 6208
rect 33134 6196 33140 6208
rect 33192 6196 33198 6248
rect 34790 6196 34796 6248
rect 34848 6236 34854 6248
rect 35253 6239 35311 6245
rect 35253 6236 35265 6239
rect 34848 6208 35265 6236
rect 34848 6196 34854 6208
rect 35253 6205 35265 6208
rect 35299 6236 35311 6239
rect 36078 6236 36084 6248
rect 35299 6208 36084 6236
rect 35299 6205 35311 6208
rect 35253 6199 35311 6205
rect 36078 6196 36084 6208
rect 36136 6196 36142 6248
rect 37829 6239 37887 6245
rect 37829 6205 37841 6239
rect 37875 6236 37887 6239
rect 37918 6236 37924 6248
rect 37875 6208 37924 6236
rect 37875 6205 37887 6208
rect 37829 6199 37887 6205
rect 37918 6196 37924 6208
rect 37976 6196 37982 6248
rect 39224 6236 39252 6276
rect 39850 6264 39856 6276
rect 39908 6264 39914 6316
rect 40402 6304 40408 6316
rect 40363 6276 40408 6304
rect 40402 6264 40408 6276
rect 40460 6264 40466 6316
rect 40512 6236 40540 6403
rect 40954 6400 40960 6412
rect 41012 6400 41018 6452
rect 41141 6443 41199 6449
rect 41141 6409 41153 6443
rect 41187 6440 41199 6443
rect 41506 6440 41512 6452
rect 41187 6412 41512 6440
rect 41187 6409 41199 6412
rect 41141 6403 41199 6409
rect 41506 6400 41512 6412
rect 41564 6400 41570 6452
rect 43898 6440 43904 6452
rect 43859 6412 43904 6440
rect 43898 6400 43904 6412
rect 43956 6400 43962 6452
rect 45002 6400 45008 6452
rect 45060 6440 45066 6452
rect 46109 6443 46167 6449
rect 46109 6440 46121 6443
rect 45060 6412 46121 6440
rect 45060 6400 45066 6412
rect 46109 6409 46121 6412
rect 46155 6409 46167 6443
rect 49878 6440 49884 6452
rect 49839 6412 49884 6440
rect 46109 6403 46167 6409
rect 49878 6400 49884 6412
rect 49936 6400 49942 6452
rect 50338 6400 50344 6452
rect 50396 6440 50402 6452
rect 51534 6440 51540 6452
rect 50396 6412 51540 6440
rect 50396 6400 50402 6412
rect 51534 6400 51540 6412
rect 51592 6400 51598 6452
rect 53282 6440 53288 6452
rect 51644 6412 53288 6440
rect 45373 6375 45431 6381
rect 45373 6341 45385 6375
rect 45419 6372 45431 6375
rect 46842 6372 46848 6384
rect 45419 6344 46848 6372
rect 45419 6341 45431 6344
rect 45373 6335 45431 6341
rect 46842 6332 46848 6344
rect 46900 6332 46906 6384
rect 47578 6332 47584 6384
rect 47636 6372 47642 6384
rect 49142 6372 49148 6384
rect 47636 6344 49148 6372
rect 47636 6332 47642 6344
rect 49142 6332 49148 6344
rect 49200 6332 49206 6384
rect 50798 6372 50804 6384
rect 50080 6344 50804 6372
rect 40589 6307 40647 6313
rect 40589 6273 40601 6307
rect 40635 6304 40647 6307
rect 41046 6304 41052 6316
rect 40635 6276 41052 6304
rect 40635 6273 40647 6276
rect 40589 6267 40647 6273
rect 41046 6264 41052 6276
rect 41104 6264 41110 6316
rect 42518 6264 42524 6316
rect 42576 6304 42582 6316
rect 42613 6307 42671 6313
rect 42613 6304 42625 6307
rect 42576 6276 42625 6304
rect 42576 6264 42582 6276
rect 42613 6273 42625 6276
rect 42659 6273 42671 6307
rect 45649 6307 45707 6313
rect 42613 6267 42671 6273
rect 42720 6276 44298 6304
rect 39224 6208 40540 6236
rect 41138 6196 41144 6248
rect 41196 6236 41202 6248
rect 42720 6236 42748 6276
rect 45649 6273 45661 6307
rect 45695 6304 45707 6307
rect 46290 6304 46296 6316
rect 45695 6276 45784 6304
rect 46251 6276 46296 6304
rect 45695 6273 45707 6276
rect 45649 6267 45707 6273
rect 41196 6208 42748 6236
rect 42889 6239 42947 6245
rect 41196 6196 41202 6208
rect 42889 6205 42901 6239
rect 42935 6236 42947 6239
rect 44910 6236 44916 6248
rect 42935 6208 44916 6236
rect 42935 6205 42947 6208
rect 42889 6199 42947 6205
rect 44910 6196 44916 6208
rect 44968 6196 44974 6248
rect 26344 6168 26372 6196
rect 28810 6168 28816 6180
rect 26344 6140 28816 6168
rect 28810 6128 28816 6140
rect 28868 6128 28874 6180
rect 35434 6128 35440 6180
rect 35492 6168 35498 6180
rect 38565 6171 38623 6177
rect 38565 6168 38577 6171
rect 35492 6140 38577 6168
rect 35492 6128 35498 6140
rect 38565 6137 38577 6140
rect 38611 6137 38623 6171
rect 38565 6131 38623 6137
rect 38654 6128 38660 6180
rect 38712 6168 38718 6180
rect 38838 6168 38844 6180
rect 38712 6140 38844 6168
rect 38712 6128 38718 6140
rect 38838 6128 38844 6140
rect 38896 6168 38902 6180
rect 41601 6171 41659 6177
rect 41601 6168 41613 6171
rect 38896 6140 41613 6168
rect 38896 6128 38902 6140
rect 41601 6137 41613 6140
rect 41647 6137 41659 6171
rect 41601 6131 41659 6137
rect 25038 6060 25044 6112
rect 25096 6100 25102 6112
rect 27890 6100 27896 6112
rect 25096 6072 27896 6100
rect 25096 6060 25102 6072
rect 27890 6060 27896 6072
rect 27948 6060 27954 6112
rect 27982 6060 27988 6112
rect 28040 6100 28046 6112
rect 28442 6100 28448 6112
rect 28040 6072 28448 6100
rect 28040 6060 28046 6072
rect 28442 6060 28448 6072
rect 28500 6060 28506 6112
rect 33962 6060 33968 6112
rect 34020 6100 34026 6112
rect 34149 6103 34207 6109
rect 34149 6100 34161 6103
rect 34020 6072 34161 6100
rect 34020 6060 34026 6072
rect 34149 6069 34161 6072
rect 34195 6100 34207 6103
rect 36170 6100 36176 6112
rect 34195 6072 36176 6100
rect 34195 6069 34207 6072
rect 34149 6063 34207 6069
rect 36170 6060 36176 6072
rect 36228 6060 36234 6112
rect 36630 6060 36636 6112
rect 36688 6100 36694 6112
rect 38010 6100 38016 6112
rect 36688 6072 38016 6100
rect 36688 6060 36694 6072
rect 38010 6060 38016 6072
rect 38068 6060 38074 6112
rect 38286 6060 38292 6112
rect 38344 6100 38350 6112
rect 39669 6103 39727 6109
rect 39669 6100 39681 6103
rect 38344 6072 39681 6100
rect 38344 6060 38350 6072
rect 39669 6069 39681 6072
rect 39715 6069 39727 6103
rect 39669 6063 39727 6069
rect 39850 6060 39856 6112
rect 39908 6100 39914 6112
rect 42610 6100 42616 6112
rect 39908 6072 42616 6100
rect 39908 6060 39914 6072
rect 42610 6060 42616 6072
rect 42668 6060 42674 6112
rect 44634 6060 44640 6112
rect 44692 6100 44698 6112
rect 45756 6100 45784 6276
rect 46290 6264 46296 6276
rect 46348 6264 46354 6316
rect 46382 6264 46388 6316
rect 46440 6304 46446 6316
rect 46569 6307 46627 6313
rect 46569 6304 46581 6307
rect 46440 6276 46581 6304
rect 46440 6264 46446 6276
rect 46569 6273 46581 6276
rect 46615 6273 46627 6307
rect 46750 6304 46756 6316
rect 46711 6276 46756 6304
rect 46569 6267 46627 6273
rect 46750 6264 46756 6276
rect 46808 6264 46814 6316
rect 47026 6264 47032 6316
rect 47084 6304 47090 6316
rect 48038 6304 48044 6316
rect 47084 6276 48044 6304
rect 47084 6264 47090 6276
rect 48038 6264 48044 6276
rect 48096 6264 48102 6316
rect 48501 6307 48559 6313
rect 48501 6273 48513 6307
rect 48547 6304 48559 6307
rect 48590 6304 48596 6316
rect 48547 6276 48596 6304
rect 48547 6273 48559 6276
rect 48501 6267 48559 6273
rect 48590 6264 48596 6276
rect 48648 6264 48654 6316
rect 50080 6313 50108 6344
rect 50798 6332 50804 6344
rect 50856 6372 50862 6384
rect 51442 6372 51448 6384
rect 50856 6344 51448 6372
rect 50856 6332 50862 6344
rect 51442 6332 51448 6344
rect 51500 6332 51506 6384
rect 49421 6307 49479 6313
rect 49421 6273 49433 6307
rect 49467 6304 49479 6307
rect 50065 6307 50123 6313
rect 49467 6276 50016 6304
rect 49467 6273 49479 6276
rect 49421 6267 49479 6273
rect 46768 6236 46796 6264
rect 49878 6236 49884 6248
rect 46768 6208 49884 6236
rect 49878 6196 49884 6208
rect 49936 6196 49942 6248
rect 47302 6128 47308 6180
rect 47360 6168 47366 6180
rect 48777 6171 48835 6177
rect 48777 6168 48789 6171
rect 47360 6140 48789 6168
rect 47360 6128 47366 6140
rect 48777 6137 48789 6140
rect 48823 6137 48835 6171
rect 48777 6131 48835 6137
rect 44692 6072 45784 6100
rect 44692 6060 44698 6072
rect 45922 6060 45928 6112
rect 45980 6100 45986 6112
rect 47857 6103 47915 6109
rect 47857 6100 47869 6103
rect 45980 6072 47869 6100
rect 45980 6060 45986 6072
rect 47857 6069 47869 6072
rect 47903 6100 47915 6103
rect 49786 6100 49792 6112
rect 47903 6072 49792 6100
rect 47903 6069 47915 6072
rect 47857 6063 47915 6069
rect 49786 6060 49792 6072
rect 49844 6060 49850 6112
rect 49988 6100 50016 6276
rect 50065 6273 50077 6307
rect 50111 6273 50123 6307
rect 50065 6267 50123 6273
rect 50154 6264 50160 6316
rect 50212 6304 50218 6316
rect 50338 6304 50344 6316
rect 50212 6276 50257 6304
rect 50299 6276 50344 6304
rect 50212 6264 50218 6276
rect 50338 6264 50344 6276
rect 50396 6264 50402 6316
rect 50525 6307 50583 6313
rect 50525 6273 50537 6307
rect 50571 6304 50583 6307
rect 50706 6304 50712 6316
rect 50571 6276 50712 6304
rect 50571 6273 50583 6276
rect 50525 6267 50583 6273
rect 50706 6264 50712 6276
rect 50764 6264 50770 6316
rect 51166 6304 51172 6316
rect 51127 6276 51172 6304
rect 51166 6264 51172 6276
rect 51224 6264 51230 6316
rect 51261 6307 51319 6313
rect 51261 6273 51273 6307
rect 51307 6304 51319 6307
rect 51644 6304 51672 6412
rect 53282 6400 53288 6412
rect 53340 6440 53346 6452
rect 54846 6440 54852 6452
rect 53340 6412 54852 6440
rect 53340 6400 53346 6412
rect 54846 6400 54852 6412
rect 54904 6440 54910 6452
rect 55033 6443 55091 6449
rect 55033 6440 55045 6443
rect 54904 6412 55045 6440
rect 54904 6400 54910 6412
rect 55033 6409 55045 6412
rect 55079 6409 55091 6443
rect 55033 6403 55091 6409
rect 58161 6443 58219 6449
rect 58161 6409 58173 6443
rect 58207 6440 58219 6443
rect 58434 6440 58440 6452
rect 58207 6412 58440 6440
rect 58207 6409 58219 6412
rect 58161 6403 58219 6409
rect 58434 6400 58440 6412
rect 58492 6400 58498 6452
rect 52178 6372 52184 6384
rect 52139 6344 52184 6372
rect 52178 6332 52184 6344
rect 52236 6332 52242 6384
rect 52270 6332 52276 6384
rect 52328 6372 52334 6384
rect 52365 6375 52423 6381
rect 52365 6372 52377 6375
rect 52328 6344 52377 6372
rect 52328 6332 52334 6344
rect 52365 6341 52377 6344
rect 52411 6341 52423 6375
rect 52365 6335 52423 6341
rect 52730 6332 52736 6384
rect 52788 6372 52794 6384
rect 54941 6375 54999 6381
rect 52788 6344 54156 6372
rect 52788 6332 52794 6344
rect 51307 6276 51672 6304
rect 51307 6273 51319 6276
rect 51261 6267 51319 6273
rect 50249 6239 50307 6245
rect 50249 6236 50261 6239
rect 50080 6208 50261 6236
rect 50080 6180 50108 6208
rect 50249 6205 50261 6208
rect 50295 6205 50307 6239
rect 50249 6199 50307 6205
rect 50430 6196 50436 6248
rect 50488 6236 50494 6248
rect 50985 6239 51043 6245
rect 50985 6236 50997 6239
rect 50488 6208 50997 6236
rect 50488 6196 50494 6208
rect 50985 6205 50997 6208
rect 51031 6205 51043 6239
rect 50985 6199 51043 6205
rect 50062 6128 50068 6180
rect 50120 6128 50126 6180
rect 51276 6168 51304 6267
rect 51718 6264 51724 6316
rect 51776 6304 51782 6316
rect 53098 6304 53104 6316
rect 51776 6276 53104 6304
rect 51776 6264 51782 6276
rect 53098 6264 53104 6276
rect 53156 6264 53162 6316
rect 54128 6313 54156 6344
rect 54941 6341 54953 6375
rect 54987 6372 54999 6375
rect 55122 6372 55128 6384
rect 54987 6344 55128 6372
rect 54987 6341 54999 6344
rect 54941 6335 54999 6341
rect 55122 6332 55128 6344
rect 55180 6332 55186 6384
rect 57514 6372 57520 6384
rect 57427 6344 57520 6372
rect 57514 6332 57520 6344
rect 57572 6372 57578 6384
rect 58342 6372 58348 6384
rect 57572 6344 58348 6372
rect 57572 6332 57578 6344
rect 58342 6332 58348 6344
rect 58400 6332 58406 6384
rect 53377 6307 53435 6313
rect 53377 6273 53389 6307
rect 53423 6273 53435 6307
rect 53377 6267 53435 6273
rect 54113 6307 54171 6313
rect 54113 6273 54125 6307
rect 54159 6273 54171 6307
rect 54113 6267 54171 6273
rect 52178 6196 52184 6248
rect 52236 6236 52242 6248
rect 52454 6236 52460 6248
rect 52236 6208 52460 6236
rect 52236 6196 52242 6208
rect 52454 6196 52460 6208
rect 52512 6196 52518 6248
rect 52914 6236 52920 6248
rect 52875 6208 52920 6236
rect 52914 6196 52920 6208
rect 52972 6196 52978 6248
rect 53006 6196 53012 6248
rect 53064 6236 53070 6248
rect 53392 6236 53420 6267
rect 54202 6236 54208 6248
rect 53064 6208 54208 6236
rect 53064 6196 53070 6208
rect 54202 6196 54208 6208
rect 54260 6196 54266 6248
rect 50264 6140 51304 6168
rect 50264 6100 50292 6140
rect 51534 6128 51540 6180
rect 51592 6168 51598 6180
rect 51997 6171 52055 6177
rect 51997 6168 52009 6171
rect 51592 6140 52009 6168
rect 51592 6128 51598 6140
rect 51997 6137 52009 6140
rect 52043 6168 52055 6171
rect 53834 6168 53840 6180
rect 52043 6140 53840 6168
rect 52043 6137 52055 6140
rect 51997 6131 52055 6137
rect 53834 6128 53840 6140
rect 53892 6128 53898 6180
rect 54297 6171 54355 6177
rect 54297 6137 54309 6171
rect 54343 6168 54355 6171
rect 56502 6168 56508 6180
rect 54343 6140 56508 6168
rect 54343 6137 54355 6140
rect 54297 6131 54355 6137
rect 56502 6128 56508 6140
rect 56560 6128 56566 6180
rect 49988 6072 50292 6100
rect 52181 6103 52239 6109
rect 52181 6069 52193 6103
rect 52227 6100 52239 6103
rect 53466 6100 53472 6112
rect 52227 6072 53472 6100
rect 52227 6069 52239 6072
rect 52181 6063 52239 6069
rect 53466 6060 53472 6072
rect 53524 6060 53530 6112
rect 54110 6060 54116 6112
rect 54168 6100 54174 6112
rect 55769 6103 55827 6109
rect 55769 6100 55781 6103
rect 54168 6072 55781 6100
rect 54168 6060 54174 6072
rect 55769 6069 55781 6072
rect 55815 6100 55827 6103
rect 56321 6103 56379 6109
rect 56321 6100 56333 6103
rect 55815 6072 56333 6100
rect 55815 6069 55827 6072
rect 55769 6063 55827 6069
rect 56321 6069 56333 6072
rect 56367 6069 56379 6103
rect 56321 6063 56379 6069
rect 56594 6060 56600 6112
rect 56652 6100 56658 6112
rect 56870 6100 56876 6112
rect 56652 6072 56876 6100
rect 56652 6060 56658 6072
rect 56870 6060 56876 6072
rect 56928 6060 56934 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 2406 5896 2412 5908
rect 2367 5868 2412 5896
rect 2406 5856 2412 5868
rect 2464 5856 2470 5908
rect 25866 5896 25872 5908
rect 25827 5868 25872 5896
rect 25866 5856 25872 5868
rect 25924 5856 25930 5908
rect 27154 5896 27160 5908
rect 27115 5868 27160 5896
rect 27154 5856 27160 5868
rect 27212 5856 27218 5908
rect 28718 5896 28724 5908
rect 28460 5868 28724 5896
rect 25774 5788 25780 5840
rect 25832 5828 25838 5840
rect 28460 5828 28488 5868
rect 28718 5856 28724 5868
rect 28776 5856 28782 5908
rect 31386 5896 31392 5908
rect 31347 5868 31392 5896
rect 31386 5856 31392 5868
rect 31444 5856 31450 5908
rect 31496 5868 31708 5896
rect 25832 5800 28488 5828
rect 25832 5788 25838 5800
rect 26513 5763 26571 5769
rect 26513 5729 26525 5763
rect 26559 5760 26571 5763
rect 27614 5760 27620 5772
rect 26559 5732 27620 5760
rect 26559 5729 26571 5732
rect 26513 5723 26571 5729
rect 27614 5720 27620 5732
rect 27672 5720 27678 5772
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2406 5692 2412 5704
rect 1903 5664 2412 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 26050 5692 26056 5704
rect 26011 5664 26056 5692
rect 26050 5652 26056 5664
rect 26108 5652 26114 5704
rect 26145 5695 26203 5701
rect 26145 5661 26157 5695
rect 26191 5692 26203 5695
rect 27338 5692 27344 5704
rect 26191 5664 26832 5692
rect 27299 5664 27344 5692
rect 26191 5661 26203 5664
rect 26145 5655 26203 5661
rect 25409 5627 25467 5633
rect 25409 5593 25421 5627
rect 25455 5624 25467 5627
rect 26160 5624 26188 5655
rect 26418 5624 26424 5636
rect 25455 5596 26188 5624
rect 26379 5596 26424 5624
rect 25455 5593 25467 5596
rect 25409 5587 25467 5593
rect 26418 5584 26424 5596
rect 26476 5584 26482 5636
rect 26804 5624 26832 5664
rect 27338 5652 27344 5664
rect 27396 5652 27402 5704
rect 27706 5692 27712 5704
rect 27667 5664 27712 5692
rect 27706 5652 27712 5664
rect 27764 5652 27770 5704
rect 28460 5701 28488 5800
rect 28626 5788 28632 5840
rect 28684 5828 28690 5840
rect 29546 5828 29552 5840
rect 28684 5800 29552 5828
rect 28684 5788 28690 5800
rect 29546 5788 29552 5800
rect 29604 5788 29610 5840
rect 30742 5788 30748 5840
rect 30800 5828 30806 5840
rect 31496 5828 31524 5868
rect 31680 5837 31708 5868
rect 32214 5856 32220 5908
rect 32272 5896 32278 5908
rect 34054 5896 34060 5908
rect 32272 5868 33640 5896
rect 34015 5868 34060 5896
rect 32272 5856 32278 5868
rect 30800 5800 31524 5828
rect 31665 5831 31723 5837
rect 30800 5788 30806 5800
rect 31665 5797 31677 5831
rect 31711 5797 31723 5831
rect 32950 5828 32956 5840
rect 31665 5791 31723 5797
rect 32048 5800 32956 5828
rect 32048 5772 32076 5800
rect 32950 5788 32956 5800
rect 33008 5788 33014 5840
rect 31757 5763 31815 5769
rect 31757 5729 31769 5763
rect 31803 5760 31815 5763
rect 32030 5760 32036 5772
rect 31803 5732 32036 5760
rect 31803 5729 31815 5732
rect 31757 5723 31815 5729
rect 32030 5720 32036 5732
rect 32088 5720 32094 5772
rect 32582 5760 32588 5772
rect 32543 5732 32588 5760
rect 32582 5720 32588 5732
rect 32640 5720 32646 5772
rect 33134 5760 33140 5772
rect 33095 5732 33140 5760
rect 33134 5720 33140 5732
rect 33192 5720 33198 5772
rect 33612 5760 33640 5868
rect 34054 5856 34060 5868
rect 34112 5856 34118 5908
rect 34422 5856 34428 5908
rect 34480 5896 34486 5908
rect 35618 5896 35624 5908
rect 34480 5868 35624 5896
rect 34480 5856 34486 5868
rect 35618 5856 35624 5868
rect 35676 5896 35682 5908
rect 37553 5899 37611 5905
rect 35676 5868 37044 5896
rect 35676 5856 35682 5868
rect 36906 5828 36912 5840
rect 36280 5800 36912 5828
rect 35158 5760 35164 5772
rect 33336 5732 33548 5760
rect 33612 5732 35164 5760
rect 27801 5695 27859 5701
rect 27801 5661 27813 5695
rect 27847 5692 27859 5695
rect 28261 5695 28319 5701
rect 28261 5692 28273 5695
rect 27847 5664 28273 5692
rect 27847 5661 27859 5664
rect 27801 5655 27859 5661
rect 28261 5661 28273 5664
rect 28307 5661 28319 5695
rect 28261 5655 28319 5661
rect 28445 5695 28503 5701
rect 28445 5661 28457 5695
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 28626 5652 28632 5704
rect 28684 5692 28690 5704
rect 28721 5695 28779 5701
rect 28721 5692 28733 5695
rect 28684 5664 28733 5692
rect 28684 5652 28690 5664
rect 28721 5661 28733 5664
rect 28767 5661 28779 5695
rect 28721 5655 28779 5661
rect 29638 5652 29644 5704
rect 29696 5692 29702 5704
rect 30009 5695 30067 5701
rect 30009 5692 30021 5695
rect 29696 5664 30021 5692
rect 29696 5652 29702 5664
rect 30009 5661 30021 5664
rect 30055 5661 30067 5695
rect 30009 5655 30067 5661
rect 30101 5695 30159 5701
rect 30101 5661 30113 5695
rect 30147 5661 30159 5695
rect 30101 5655 30159 5661
rect 28534 5624 28540 5636
rect 26804 5596 28540 5624
rect 28534 5584 28540 5596
rect 28592 5584 28598 5636
rect 30116 5624 30144 5655
rect 30190 5652 30196 5704
rect 30248 5692 30254 5704
rect 30377 5695 30435 5701
rect 30248 5664 30293 5692
rect 30248 5652 30254 5664
rect 30377 5661 30389 5695
rect 30423 5692 30435 5695
rect 30558 5692 30564 5704
rect 30423 5664 30564 5692
rect 30423 5661 30435 5664
rect 30377 5655 30435 5661
rect 30558 5652 30564 5664
rect 30616 5652 30622 5704
rect 31573 5695 31631 5701
rect 31573 5661 31585 5695
rect 31619 5661 31631 5695
rect 31573 5655 31631 5661
rect 31588 5624 31616 5655
rect 31846 5652 31852 5704
rect 31904 5692 31910 5704
rect 33336 5701 33364 5732
rect 33321 5695 33379 5701
rect 31904 5664 31949 5692
rect 31904 5652 31910 5664
rect 33321 5661 33333 5695
rect 33367 5661 33379 5695
rect 33321 5655 33379 5661
rect 33413 5695 33471 5701
rect 33413 5661 33425 5695
rect 33459 5661 33471 5695
rect 33413 5655 33471 5661
rect 33042 5624 33048 5636
rect 28966 5596 33048 5624
rect 28966 5590 28994 5596
rect 28736 5568 28994 5590
rect 33042 5584 33048 5596
rect 33100 5584 33106 5636
rect 33226 5584 33232 5636
rect 33284 5624 33290 5636
rect 33428 5624 33456 5655
rect 33284 5596 33456 5624
rect 33520 5624 33548 5732
rect 35158 5720 35164 5732
rect 35216 5720 35222 5772
rect 35342 5760 35348 5772
rect 35268 5732 35348 5760
rect 34238 5652 34244 5704
rect 34296 5692 34302 5704
rect 35268 5701 35296 5732
rect 35342 5720 35348 5732
rect 35400 5760 35406 5772
rect 36280 5769 36308 5800
rect 36906 5788 36912 5800
rect 36964 5788 36970 5840
rect 37016 5828 37044 5868
rect 37553 5865 37565 5899
rect 37599 5896 37611 5899
rect 39482 5896 39488 5908
rect 37599 5868 39488 5896
rect 37599 5865 37611 5868
rect 37553 5859 37611 5865
rect 39482 5856 39488 5868
rect 39540 5856 39546 5908
rect 42150 5896 42156 5908
rect 42111 5868 42156 5896
rect 42150 5856 42156 5868
rect 42208 5896 42214 5908
rect 42794 5896 42800 5908
rect 42208 5868 42800 5896
rect 42208 5856 42214 5868
rect 42794 5856 42800 5868
rect 42852 5856 42858 5908
rect 46198 5856 46204 5908
rect 46256 5896 46262 5908
rect 46753 5899 46811 5905
rect 46753 5896 46765 5899
rect 46256 5868 46765 5896
rect 46256 5856 46262 5868
rect 46753 5865 46765 5868
rect 46799 5865 46811 5899
rect 48774 5896 48780 5908
rect 46753 5859 46811 5865
rect 47044 5868 48780 5896
rect 40678 5828 40684 5840
rect 37016 5800 40684 5828
rect 40678 5788 40684 5800
rect 40736 5788 40742 5840
rect 41414 5788 41420 5840
rect 41472 5828 41478 5840
rect 44269 5831 44327 5837
rect 41472 5800 41644 5828
rect 41472 5788 41478 5800
rect 36265 5763 36323 5769
rect 36265 5760 36277 5763
rect 35400 5732 36277 5760
rect 35400 5720 35406 5732
rect 36265 5729 36277 5732
rect 36311 5729 36323 5763
rect 36265 5723 36323 5729
rect 36354 5720 36360 5772
rect 36412 5760 36418 5772
rect 36998 5760 37004 5772
rect 36412 5732 36457 5760
rect 36959 5732 37004 5760
rect 36412 5720 36418 5732
rect 36998 5720 37004 5732
rect 37056 5720 37062 5772
rect 41616 5769 41644 5800
rect 44269 5797 44281 5831
rect 44315 5828 44327 5831
rect 45373 5831 45431 5837
rect 45373 5828 45385 5831
rect 44315 5800 45385 5828
rect 44315 5797 44327 5800
rect 44269 5791 44327 5797
rect 45373 5797 45385 5800
rect 45419 5797 45431 5831
rect 45373 5791 45431 5797
rect 37093 5763 37151 5769
rect 37093 5729 37105 5763
rect 37139 5760 37151 5763
rect 41233 5763 41291 5769
rect 37139 5732 38516 5760
rect 37139 5729 37151 5732
rect 37093 5723 37151 5729
rect 38488 5704 38516 5732
rect 41233 5729 41245 5763
rect 41279 5760 41291 5763
rect 41601 5763 41659 5769
rect 41279 5732 41460 5760
rect 41279 5729 41291 5732
rect 41233 5723 41291 5729
rect 35253 5695 35311 5701
rect 35253 5692 35265 5695
rect 34296 5664 35265 5692
rect 34296 5652 34302 5664
rect 35253 5661 35265 5664
rect 35299 5661 35311 5695
rect 35253 5655 35311 5661
rect 35955 5695 36013 5701
rect 35955 5661 35967 5695
rect 36001 5692 36013 5695
rect 36170 5692 36176 5704
rect 36001 5664 36176 5692
rect 36001 5661 36013 5664
rect 35955 5655 36013 5661
rect 36170 5652 36176 5664
rect 36228 5652 36234 5704
rect 38010 5692 38016 5704
rect 37971 5664 38016 5692
rect 38010 5652 38016 5664
rect 38068 5652 38074 5704
rect 38194 5701 38200 5704
rect 38171 5695 38200 5701
rect 38171 5661 38183 5695
rect 38171 5655 38200 5661
rect 38186 5652 38200 5655
rect 38252 5652 38258 5704
rect 38286 5652 38292 5704
rect 38344 5692 38350 5704
rect 38344 5664 38389 5692
rect 38344 5652 38350 5664
rect 38470 5652 38476 5704
rect 38528 5692 38534 5704
rect 39114 5692 39120 5704
rect 38528 5664 39120 5692
rect 38528 5652 38534 5664
rect 39114 5652 39120 5664
rect 39172 5652 39178 5704
rect 39301 5695 39359 5701
rect 39301 5661 39313 5695
rect 39347 5692 39359 5695
rect 39390 5692 39396 5704
rect 39347 5664 39396 5692
rect 39347 5661 39359 5664
rect 39301 5655 39359 5661
rect 39390 5652 39396 5664
rect 39448 5652 39454 5704
rect 40034 5652 40040 5704
rect 40092 5692 40098 5704
rect 41138 5692 41144 5704
rect 40092 5664 41144 5692
rect 40092 5652 40098 5664
rect 41138 5652 41144 5664
rect 41196 5652 41202 5704
rect 41322 5692 41328 5704
rect 41283 5664 41328 5692
rect 41322 5652 41328 5664
rect 41380 5652 41386 5704
rect 34606 5624 34612 5636
rect 33520 5596 34612 5624
rect 33284 5584 33290 5596
rect 34606 5584 34612 5596
rect 34664 5584 34670 5636
rect 36998 5624 37004 5636
rect 35452 5596 37004 5624
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 27338 5556 27344 5568
rect 27299 5528 27344 5556
rect 27338 5516 27344 5528
rect 27396 5516 27402 5568
rect 28350 5516 28356 5568
rect 28408 5556 28414 5568
rect 28629 5559 28687 5565
rect 28629 5556 28641 5559
rect 28408 5528 28641 5556
rect 28408 5516 28414 5528
rect 28629 5525 28641 5528
rect 28675 5525 28687 5559
rect 28629 5519 28687 5525
rect 28718 5516 28724 5568
rect 28776 5562 28994 5568
rect 28776 5516 28782 5562
rect 29546 5516 29552 5568
rect 29604 5556 29610 5568
rect 29733 5559 29791 5565
rect 29733 5556 29745 5559
rect 29604 5528 29745 5556
rect 29604 5516 29610 5528
rect 29733 5525 29745 5528
rect 29779 5525 29791 5559
rect 29733 5519 29791 5525
rect 34698 5516 34704 5568
rect 34756 5556 34762 5568
rect 35066 5556 35072 5568
rect 34756 5528 35072 5556
rect 34756 5516 34762 5528
rect 35066 5516 35072 5528
rect 35124 5516 35130 5568
rect 35250 5516 35256 5568
rect 35308 5556 35314 5568
rect 35452 5556 35480 5596
rect 36998 5584 37004 5596
rect 37056 5584 37062 5636
rect 37185 5627 37243 5633
rect 37185 5593 37197 5627
rect 37231 5624 37243 5627
rect 38186 5624 38214 5652
rect 37231 5596 38214 5624
rect 38381 5627 38439 5633
rect 37231 5593 37243 5596
rect 37185 5587 37243 5593
rect 38381 5593 38393 5627
rect 38427 5624 38439 5627
rect 39209 5627 39267 5633
rect 39209 5624 39221 5627
rect 38427 5596 39221 5624
rect 38427 5593 38439 5596
rect 38381 5587 38439 5593
rect 39209 5593 39221 5596
rect 39255 5593 39267 5627
rect 41230 5624 41236 5636
rect 39209 5587 39267 5593
rect 39960 5596 41236 5624
rect 35308 5528 35480 5556
rect 35308 5516 35314 5528
rect 35710 5516 35716 5568
rect 35768 5556 35774 5568
rect 35805 5559 35863 5565
rect 35805 5556 35817 5559
rect 35768 5528 35817 5556
rect 35768 5516 35774 5528
rect 35805 5525 35817 5528
rect 35851 5525 35863 5559
rect 35805 5519 35863 5525
rect 38657 5559 38715 5565
rect 38657 5525 38669 5559
rect 38703 5556 38715 5559
rect 39960 5556 39988 5596
rect 41230 5584 41236 5596
rect 41288 5584 41294 5636
rect 41432 5624 41460 5732
rect 41601 5729 41613 5763
rect 41647 5729 41659 5763
rect 41601 5723 41659 5729
rect 41693 5763 41751 5769
rect 41693 5729 41705 5763
rect 41739 5760 41751 5763
rect 43162 5760 43168 5772
rect 41739 5732 43168 5760
rect 41739 5729 41751 5732
rect 41693 5723 41751 5729
rect 43162 5720 43168 5732
rect 43220 5720 43226 5772
rect 43346 5760 43352 5772
rect 43307 5732 43352 5760
rect 43346 5720 43352 5732
rect 43404 5720 43410 5772
rect 45278 5760 45284 5772
rect 45239 5732 45284 5760
rect 45278 5720 45284 5732
rect 45336 5760 45342 5772
rect 46382 5760 46388 5772
rect 45336 5732 46388 5760
rect 45336 5720 45342 5732
rect 46382 5720 46388 5732
rect 46440 5720 46446 5772
rect 47044 5760 47072 5868
rect 48774 5856 48780 5868
rect 48832 5896 48838 5908
rect 50430 5896 50436 5908
rect 48832 5868 50436 5896
rect 48832 5856 48838 5868
rect 50430 5856 50436 5868
rect 50488 5856 50494 5908
rect 50525 5899 50583 5905
rect 50525 5865 50537 5899
rect 50571 5896 50583 5899
rect 50982 5896 50988 5908
rect 50571 5868 50988 5896
rect 50571 5865 50583 5868
rect 50525 5859 50583 5865
rect 50982 5856 50988 5868
rect 51040 5856 51046 5908
rect 51537 5899 51595 5905
rect 51537 5865 51549 5899
rect 51583 5896 51595 5899
rect 52362 5896 52368 5908
rect 51583 5868 52368 5896
rect 51583 5865 51595 5868
rect 51537 5859 51595 5865
rect 48314 5828 48320 5840
rect 48275 5800 48320 5828
rect 48314 5788 48320 5800
rect 48372 5788 48378 5840
rect 50614 5828 50620 5840
rect 50575 5800 50620 5828
rect 50614 5788 50620 5800
rect 50672 5788 50678 5840
rect 51552 5828 51580 5859
rect 52362 5856 52368 5868
rect 52420 5856 52426 5908
rect 52914 5856 52920 5908
rect 52972 5896 52978 5908
rect 53558 5896 53564 5908
rect 52972 5868 53564 5896
rect 52972 5856 52978 5868
rect 53558 5856 53564 5868
rect 53616 5896 53622 5908
rect 56045 5899 56103 5905
rect 56045 5896 56057 5899
rect 53616 5868 56057 5896
rect 53616 5856 53622 5868
rect 56045 5865 56057 5868
rect 56091 5865 56103 5899
rect 56045 5859 56103 5865
rect 56502 5856 56508 5908
rect 56560 5896 56566 5908
rect 56597 5899 56655 5905
rect 56597 5896 56609 5899
rect 56560 5868 56609 5896
rect 56560 5856 56566 5868
rect 56597 5865 56609 5868
rect 56643 5865 56655 5899
rect 57146 5896 57152 5908
rect 57107 5868 57152 5896
rect 56597 5859 56655 5865
rect 57146 5856 57152 5868
rect 57204 5856 57210 5908
rect 58345 5899 58403 5905
rect 58345 5865 58357 5899
rect 58391 5896 58403 5899
rect 58526 5896 58532 5908
rect 58391 5868 58532 5896
rect 58391 5865 58403 5868
rect 58345 5859 58403 5865
rect 58526 5856 58532 5868
rect 58584 5856 58590 5908
rect 55490 5828 55496 5840
rect 50724 5800 51580 5828
rect 55451 5800 55496 5828
rect 48685 5763 48743 5769
rect 46952 5732 47072 5760
rect 47320 5732 48314 5760
rect 43254 5692 43260 5704
rect 43215 5664 43260 5692
rect 43254 5652 43260 5664
rect 43312 5652 43318 5704
rect 43364 5692 43392 5720
rect 43993 5695 44051 5701
rect 43993 5692 44005 5695
rect 43364 5664 44005 5692
rect 43993 5661 44005 5664
rect 44039 5661 44051 5695
rect 45189 5695 45247 5701
rect 45189 5692 45201 5695
rect 43993 5655 44051 5661
rect 44100 5664 45201 5692
rect 42058 5624 42064 5636
rect 41432 5596 42064 5624
rect 42058 5584 42064 5596
rect 42116 5584 42122 5636
rect 42978 5584 42984 5636
rect 43036 5624 43042 5636
rect 44100 5624 44128 5664
rect 45189 5661 45201 5664
rect 45235 5661 45247 5695
rect 45462 5692 45468 5704
rect 45189 5655 45247 5661
rect 45388 5664 45468 5692
rect 44266 5624 44272 5636
rect 43036 5596 44128 5624
rect 44227 5596 44272 5624
rect 43036 5584 43042 5596
rect 44266 5584 44272 5596
rect 44324 5584 44330 5636
rect 44910 5584 44916 5636
rect 44968 5624 44974 5636
rect 45388 5624 45416 5664
rect 45462 5652 45468 5664
rect 45520 5652 45526 5704
rect 46952 5701 46980 5732
rect 46937 5695 46995 5701
rect 45572 5664 46888 5692
rect 45572 5624 45600 5664
rect 44968 5596 45416 5624
rect 45480 5596 45600 5624
rect 44968 5584 44974 5596
rect 38703 5528 39988 5556
rect 40129 5559 40187 5565
rect 38703 5525 38715 5528
rect 38657 5519 38715 5525
rect 40129 5525 40141 5559
rect 40175 5556 40187 5559
rect 40678 5556 40684 5568
rect 40175 5528 40684 5556
rect 40175 5525 40187 5528
rect 40129 5519 40187 5525
rect 40678 5516 40684 5528
rect 40736 5516 40742 5568
rect 41046 5556 41052 5568
rect 41007 5528 41052 5556
rect 41046 5516 41052 5528
rect 41104 5516 41110 5568
rect 42334 5516 42340 5568
rect 42392 5556 42398 5568
rect 42889 5559 42947 5565
rect 42889 5556 42901 5559
rect 42392 5528 42901 5556
rect 42392 5516 42398 5528
rect 42889 5525 42901 5528
rect 42935 5525 42947 5559
rect 42889 5519 42947 5525
rect 43990 5516 43996 5568
rect 44048 5556 44054 5568
rect 44085 5559 44143 5565
rect 44085 5556 44097 5559
rect 44048 5528 44097 5556
rect 44048 5516 44054 5528
rect 44085 5525 44097 5528
rect 44131 5556 44143 5559
rect 45480 5556 45508 5596
rect 45646 5584 45652 5636
rect 45704 5624 45710 5636
rect 46860 5624 46888 5664
rect 46937 5661 46949 5695
rect 46983 5661 46995 5695
rect 46937 5655 46995 5661
rect 47029 5695 47087 5701
rect 47029 5661 47041 5695
rect 47075 5692 47087 5695
rect 47210 5692 47216 5704
rect 47075 5664 47216 5692
rect 47075 5661 47087 5664
rect 47029 5655 47087 5661
rect 47210 5652 47216 5664
rect 47268 5652 47274 5704
rect 47320 5701 47348 5732
rect 47305 5695 47363 5701
rect 47305 5661 47317 5695
rect 47351 5661 47363 5695
rect 47305 5655 47363 5661
rect 47397 5695 47455 5701
rect 47397 5661 47409 5695
rect 47443 5692 47455 5695
rect 47762 5692 47768 5704
rect 47443 5664 47768 5692
rect 47443 5661 47455 5664
rect 47397 5655 47455 5661
rect 47762 5652 47768 5664
rect 47820 5652 47826 5704
rect 48038 5692 48044 5704
rect 47999 5664 48044 5692
rect 48038 5652 48044 5664
rect 48096 5652 48102 5704
rect 47121 5627 47179 5633
rect 45704 5596 45749 5624
rect 46860 5596 46980 5624
rect 45704 5584 45710 5596
rect 46952 5568 46980 5596
rect 47121 5593 47133 5627
rect 47167 5624 47179 5627
rect 47486 5624 47492 5636
rect 47167 5596 47492 5624
rect 47167 5593 47179 5596
rect 47121 5587 47179 5593
rect 47486 5584 47492 5596
rect 47544 5584 47550 5636
rect 48286 5624 48314 5732
rect 48685 5729 48697 5763
rect 48731 5760 48743 5763
rect 48774 5760 48780 5772
rect 48731 5732 48780 5760
rect 48731 5729 48743 5732
rect 48685 5723 48743 5729
rect 48774 5720 48780 5732
rect 48832 5720 48838 5772
rect 49878 5720 49884 5772
rect 49936 5760 49942 5772
rect 50724 5760 50752 5800
rect 55490 5788 55496 5800
rect 55548 5788 55554 5840
rect 49936 5732 50752 5760
rect 49936 5720 49942 5732
rect 51902 5720 51908 5772
rect 51960 5760 51966 5772
rect 52181 5763 52239 5769
rect 52181 5760 52193 5763
rect 51960 5732 52193 5760
rect 51960 5720 51966 5732
rect 52181 5729 52193 5732
rect 52227 5729 52239 5763
rect 53098 5760 53104 5772
rect 53059 5732 53104 5760
rect 52181 5723 52239 5729
rect 53098 5720 53104 5732
rect 53156 5720 53162 5772
rect 54110 5760 54116 5772
rect 54023 5732 54116 5760
rect 54110 5720 54116 5732
rect 54168 5760 54174 5772
rect 54754 5760 54760 5772
rect 54168 5732 54760 5760
rect 54168 5720 54174 5732
rect 54754 5720 54760 5732
rect 54812 5720 54818 5772
rect 55030 5720 55036 5772
rect 55088 5760 55094 5772
rect 57701 5763 57759 5769
rect 57701 5760 57713 5763
rect 55088 5732 57713 5760
rect 55088 5720 55094 5732
rect 57701 5729 57713 5732
rect 57747 5729 57759 5763
rect 57701 5723 57759 5729
rect 48590 5692 48596 5704
rect 48551 5664 48596 5692
rect 48590 5652 48596 5664
rect 48648 5652 48654 5704
rect 49329 5695 49387 5701
rect 49329 5661 49341 5695
rect 49375 5692 49387 5695
rect 49602 5692 49608 5704
rect 49375 5664 49608 5692
rect 49375 5661 49387 5664
rect 49329 5655 49387 5661
rect 49602 5652 49608 5664
rect 49660 5652 49666 5704
rect 50890 5652 50896 5704
rect 50948 5692 50954 5704
rect 50985 5695 51043 5701
rect 50985 5692 50997 5695
rect 50948 5664 50997 5692
rect 50948 5652 50954 5664
rect 50985 5661 50997 5664
rect 51031 5692 51043 5695
rect 52457 5695 52515 5701
rect 52457 5692 52469 5695
rect 51031 5664 52469 5692
rect 51031 5661 51043 5664
rect 50985 5655 51043 5661
rect 52457 5661 52469 5664
rect 52503 5661 52515 5695
rect 52457 5655 52515 5661
rect 53377 5695 53435 5701
rect 53377 5661 53389 5695
rect 53423 5692 53435 5695
rect 53466 5692 53472 5704
rect 53423 5664 53472 5692
rect 53423 5661 53435 5664
rect 53377 5655 53435 5661
rect 48682 5624 48688 5636
rect 48286 5596 48688 5624
rect 48682 5584 48688 5596
rect 48740 5584 48746 5636
rect 52472 5624 52500 5655
rect 53466 5652 53472 5664
rect 53524 5652 53530 5704
rect 54202 5692 54208 5704
rect 54163 5664 54208 5692
rect 54202 5652 54208 5664
rect 54260 5652 54266 5704
rect 54846 5692 54852 5704
rect 54807 5664 54852 5692
rect 54846 5652 54852 5664
rect 54904 5652 54910 5704
rect 55122 5624 55128 5636
rect 52472 5596 55128 5624
rect 55122 5584 55128 5596
rect 55180 5584 55186 5636
rect 44131 5528 45508 5556
rect 45557 5559 45615 5565
rect 44131 5525 44143 5528
rect 44085 5519 44143 5525
rect 45557 5525 45569 5559
rect 45603 5556 45615 5559
rect 45738 5556 45744 5568
rect 45603 5528 45744 5556
rect 45603 5525 45615 5528
rect 45557 5519 45615 5525
rect 45738 5516 45744 5528
rect 45796 5556 45802 5568
rect 46014 5556 46020 5568
rect 45796 5528 46020 5556
rect 45796 5516 45802 5528
rect 46014 5516 46020 5528
rect 46072 5556 46078 5568
rect 46109 5559 46167 5565
rect 46109 5556 46121 5559
rect 46072 5528 46121 5556
rect 46072 5516 46078 5528
rect 46109 5525 46121 5528
rect 46155 5525 46167 5559
rect 46109 5519 46167 5525
rect 46934 5516 46940 5568
rect 46992 5516 46998 5568
rect 48700 5556 48728 5584
rect 52914 5556 52920 5568
rect 48700 5528 52920 5556
rect 52914 5516 52920 5528
rect 52972 5516 52978 5568
rect 54846 5556 54852 5568
rect 54807 5528 54852 5556
rect 54846 5516 54852 5528
rect 54904 5516 54910 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 26142 5352 26148 5364
rect 26103 5324 26148 5352
rect 26142 5312 26148 5324
rect 26200 5312 26206 5364
rect 27338 5352 27344 5364
rect 27299 5324 27344 5352
rect 27338 5312 27344 5324
rect 27396 5312 27402 5364
rect 28810 5352 28816 5364
rect 27448 5324 28816 5352
rect 25958 5244 25964 5296
rect 26016 5284 26022 5296
rect 27448 5284 27476 5324
rect 28810 5312 28816 5324
rect 28868 5352 28874 5364
rect 28921 5355 28979 5361
rect 28921 5352 28933 5355
rect 28868 5324 28933 5352
rect 28868 5312 28874 5324
rect 28921 5321 28933 5324
rect 28967 5321 28979 5355
rect 28921 5315 28979 5321
rect 29089 5355 29147 5361
rect 29089 5321 29101 5355
rect 29135 5321 29147 5355
rect 30098 5352 30104 5364
rect 30059 5324 30104 5352
rect 29089 5315 29147 5321
rect 26016 5256 27476 5284
rect 28721 5287 28779 5293
rect 26016 5244 26022 5256
rect 28721 5253 28733 5287
rect 28767 5253 28779 5287
rect 29104 5284 29132 5315
rect 30098 5312 30104 5324
rect 30156 5312 30162 5364
rect 31757 5355 31815 5361
rect 31757 5321 31769 5355
rect 31803 5352 31815 5355
rect 31846 5352 31852 5364
rect 31803 5324 31852 5352
rect 31803 5321 31815 5324
rect 31757 5315 31815 5321
rect 31846 5312 31852 5324
rect 31904 5312 31910 5364
rect 32769 5355 32827 5361
rect 32769 5321 32781 5355
rect 32815 5352 32827 5355
rect 33042 5352 33048 5364
rect 32815 5324 33048 5352
rect 32815 5321 32827 5324
rect 32769 5315 32827 5321
rect 33042 5312 33048 5324
rect 33100 5312 33106 5364
rect 33778 5352 33784 5364
rect 33739 5324 33784 5352
rect 33778 5312 33784 5324
rect 33836 5352 33842 5364
rect 36265 5355 36323 5361
rect 33836 5324 36232 5352
rect 33836 5312 33842 5324
rect 29104 5256 29684 5284
rect 28721 5247 28779 5253
rect 26326 5176 26332 5228
rect 26384 5216 26390 5228
rect 26421 5219 26479 5225
rect 26421 5216 26433 5219
rect 26384 5188 26433 5216
rect 26384 5176 26390 5188
rect 26421 5185 26433 5188
rect 26467 5185 26479 5219
rect 26421 5179 26479 5185
rect 26786 5176 26792 5228
rect 26844 5216 26850 5228
rect 27433 5219 27491 5225
rect 27433 5216 27445 5219
rect 26844 5188 27445 5216
rect 26844 5176 26850 5188
rect 27433 5185 27445 5188
rect 27479 5185 27491 5219
rect 27433 5179 27491 5185
rect 27617 5219 27675 5225
rect 27617 5185 27629 5219
rect 27663 5185 27675 5219
rect 27798 5216 27804 5228
rect 27759 5188 27804 5216
rect 27617 5179 27675 5185
rect 26970 5108 26976 5160
rect 27028 5148 27034 5160
rect 27341 5151 27399 5157
rect 27341 5148 27353 5151
rect 27028 5120 27353 5148
rect 27028 5108 27034 5120
rect 27341 5117 27353 5120
rect 27387 5117 27399 5151
rect 27632 5148 27660 5179
rect 27798 5176 27804 5188
rect 27856 5176 27862 5228
rect 28736 5216 28764 5247
rect 29362 5216 29368 5228
rect 28736 5188 29368 5216
rect 29362 5176 29368 5188
rect 29420 5176 29426 5228
rect 29546 5216 29552 5228
rect 29507 5188 29552 5216
rect 29546 5176 29552 5188
rect 29604 5176 29610 5228
rect 29656 5225 29684 5256
rect 30190 5244 30196 5296
rect 30248 5284 30254 5296
rect 32306 5284 32312 5296
rect 30248 5256 32312 5284
rect 30248 5244 30254 5256
rect 29641 5219 29699 5225
rect 29641 5185 29653 5219
rect 29687 5185 29699 5219
rect 29641 5179 29699 5185
rect 29825 5219 29883 5225
rect 29825 5185 29837 5219
rect 29871 5185 29883 5219
rect 29825 5179 29883 5185
rect 29917 5219 29975 5225
rect 29917 5185 29929 5219
rect 29963 5216 29975 5219
rect 30742 5216 30748 5228
rect 29963 5188 30748 5216
rect 29963 5185 29975 5188
rect 29917 5179 29975 5185
rect 29178 5148 29184 5160
rect 27632 5120 29184 5148
rect 27341 5111 27399 5117
rect 29178 5108 29184 5120
rect 29236 5108 29242 5160
rect 29840 5148 29868 5179
rect 30742 5176 30748 5188
rect 30800 5176 30806 5228
rect 31113 5219 31171 5225
rect 31113 5185 31125 5219
rect 31159 5185 31171 5219
rect 31294 5216 31300 5228
rect 31255 5188 31300 5216
rect 31113 5179 31171 5185
rect 31128 5148 31156 5179
rect 31294 5176 31300 5188
rect 31352 5176 31358 5228
rect 31404 5225 31432 5256
rect 32306 5244 32312 5256
rect 32364 5284 32370 5296
rect 32490 5284 32496 5296
rect 32364 5256 32496 5284
rect 32364 5244 32370 5256
rect 32490 5244 32496 5256
rect 32548 5244 32554 5296
rect 35802 5244 35808 5296
rect 35860 5244 35866 5296
rect 31389 5219 31447 5225
rect 31389 5185 31401 5219
rect 31435 5185 31447 5219
rect 31389 5179 31447 5185
rect 31478 5176 31484 5228
rect 31536 5216 31542 5228
rect 31846 5216 31852 5228
rect 31536 5188 31852 5216
rect 31536 5176 31542 5188
rect 31846 5176 31852 5188
rect 31904 5176 31910 5228
rect 32674 5216 32680 5228
rect 31956 5188 32680 5216
rect 31956 5148 31984 5188
rect 32674 5176 32680 5188
rect 32732 5176 32738 5228
rect 33689 5219 33747 5225
rect 33689 5216 33701 5219
rect 33152 5188 33701 5216
rect 33152 5148 33180 5188
rect 33689 5185 33701 5188
rect 33735 5185 33747 5219
rect 33689 5179 33747 5185
rect 33873 5219 33931 5225
rect 33873 5185 33885 5219
rect 33919 5185 33931 5219
rect 36204 5216 36232 5324
rect 36265 5321 36277 5355
rect 36311 5352 36323 5355
rect 41417 5355 41475 5361
rect 41417 5352 41429 5355
rect 36311 5324 41429 5352
rect 36311 5321 36323 5324
rect 36265 5315 36323 5321
rect 41417 5321 41429 5324
rect 41463 5321 41475 5355
rect 45649 5355 45707 5361
rect 45649 5352 45661 5355
rect 41417 5315 41475 5321
rect 43088 5324 45661 5352
rect 36817 5287 36875 5293
rect 36817 5253 36829 5287
rect 36863 5284 36875 5287
rect 37642 5284 37648 5296
rect 36863 5256 37648 5284
rect 36863 5253 36875 5256
rect 36817 5247 36875 5253
rect 37642 5244 37648 5256
rect 37700 5244 37706 5296
rect 38194 5284 38200 5296
rect 37752 5256 38200 5284
rect 37752 5225 37780 5256
rect 38194 5244 38200 5256
rect 38252 5244 38258 5296
rect 40034 5284 40040 5296
rect 39882 5256 40040 5284
rect 40034 5244 40040 5256
rect 40092 5244 40098 5296
rect 40313 5287 40371 5293
rect 40313 5253 40325 5287
rect 40359 5284 40371 5287
rect 41046 5284 41052 5296
rect 40359 5256 41052 5284
rect 40359 5253 40371 5256
rect 40313 5247 40371 5253
rect 41046 5244 41052 5256
rect 41104 5244 41110 5296
rect 41432 5284 41460 5315
rect 41782 5284 41788 5296
rect 41432 5256 41788 5284
rect 41782 5244 41788 5256
rect 41840 5244 41846 5296
rect 42613 5287 42671 5293
rect 42613 5253 42625 5287
rect 42659 5284 42671 5287
rect 42794 5284 42800 5296
rect 42659 5256 42800 5284
rect 42659 5253 42671 5256
rect 42613 5247 42671 5253
rect 42794 5244 42800 5256
rect 42852 5244 42858 5296
rect 37737 5219 37795 5225
rect 36204 5188 37320 5216
rect 33873 5179 33931 5185
rect 29840 5120 31984 5148
rect 32048 5120 33180 5148
rect 27525 5083 27583 5089
rect 27525 5049 27537 5083
rect 27571 5080 27583 5083
rect 27982 5080 27988 5092
rect 27571 5052 27988 5080
rect 27571 5049 27583 5052
rect 27525 5043 27583 5049
rect 27982 5040 27988 5052
rect 28040 5040 28046 5092
rect 28258 5040 28264 5092
rect 28316 5080 28322 5092
rect 30466 5080 30472 5092
rect 28316 5052 30472 5080
rect 28316 5040 28322 5052
rect 30466 5040 30472 5052
rect 30524 5080 30530 5092
rect 32048 5080 32076 5120
rect 33226 5108 33232 5160
rect 33284 5148 33290 5160
rect 33284 5120 33377 5148
rect 33284 5108 33290 5120
rect 33410 5108 33416 5160
rect 33468 5148 33474 5160
rect 33888 5148 33916 5179
rect 34514 5148 34520 5160
rect 33468 5120 33916 5148
rect 34475 5120 34520 5148
rect 33468 5108 33474 5120
rect 34514 5108 34520 5120
rect 34572 5108 34578 5160
rect 34793 5151 34851 5157
rect 34793 5117 34805 5151
rect 34839 5148 34851 5151
rect 37182 5148 37188 5160
rect 34839 5120 37188 5148
rect 34839 5117 34851 5120
rect 34793 5111 34851 5117
rect 37182 5108 37188 5120
rect 37240 5108 37246 5160
rect 30524 5052 32076 5080
rect 30524 5040 30530 5052
rect 32766 5040 32772 5092
rect 32824 5080 32830 5092
rect 32861 5083 32919 5089
rect 32861 5080 32873 5083
rect 32824 5052 32873 5080
rect 32824 5040 32830 5052
rect 32861 5049 32873 5052
rect 32907 5049 32919 5083
rect 32861 5043 32919 5049
rect 26878 4972 26884 5024
rect 26936 5012 26942 5024
rect 28902 5012 28908 5024
rect 26936 4984 28908 5012
rect 26936 4972 26942 4984
rect 28902 4972 28908 4984
rect 28960 4972 28966 5024
rect 30190 4972 30196 5024
rect 30248 5012 30254 5024
rect 30561 5015 30619 5021
rect 30561 5012 30573 5015
rect 30248 4984 30573 5012
rect 30248 4972 30254 4984
rect 30561 4981 30573 4984
rect 30607 4981 30619 5015
rect 30561 4975 30619 4981
rect 32306 4972 32312 5024
rect 32364 5012 32370 5024
rect 33244 5012 33272 5108
rect 37292 5080 37320 5188
rect 37737 5185 37749 5219
rect 37783 5185 37795 5219
rect 37737 5179 37795 5185
rect 37829 5219 37887 5225
rect 37829 5185 37841 5219
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 37844 5148 37872 5179
rect 37918 5176 37924 5228
rect 37976 5216 37982 5228
rect 38105 5219 38163 5225
rect 37976 5188 38021 5216
rect 37976 5176 37982 5188
rect 38105 5185 38117 5219
rect 38151 5216 38163 5219
rect 38470 5216 38476 5228
rect 38151 5188 38476 5216
rect 38151 5185 38163 5188
rect 38105 5179 38163 5185
rect 38470 5176 38476 5188
rect 38528 5176 38534 5228
rect 41414 5176 41420 5228
rect 41472 5216 41478 5228
rect 41509 5219 41567 5225
rect 41509 5216 41521 5219
rect 41472 5188 41521 5216
rect 41472 5176 41478 5188
rect 41509 5185 41521 5188
rect 41555 5216 41567 5219
rect 43088 5216 43116 5324
rect 45649 5321 45661 5324
rect 45695 5352 45707 5355
rect 46658 5352 46664 5364
rect 45695 5324 46664 5352
rect 45695 5321 45707 5324
rect 45649 5315 45707 5321
rect 46658 5312 46664 5324
rect 46716 5312 46722 5364
rect 46842 5352 46848 5364
rect 46803 5324 46848 5352
rect 46842 5312 46848 5324
rect 46900 5312 46906 5364
rect 47486 5312 47492 5364
rect 47544 5352 47550 5364
rect 48409 5355 48467 5361
rect 48409 5352 48421 5355
rect 47544 5324 48421 5352
rect 47544 5312 47550 5324
rect 48409 5321 48421 5324
rect 48455 5321 48467 5355
rect 48409 5315 48467 5321
rect 49694 5312 49700 5364
rect 49752 5352 49758 5364
rect 50249 5355 50307 5361
rect 50249 5352 50261 5355
rect 49752 5324 50261 5352
rect 49752 5312 49758 5324
rect 50249 5321 50261 5324
rect 50295 5321 50307 5355
rect 50249 5315 50307 5321
rect 50798 5312 50804 5364
rect 50856 5352 50862 5364
rect 51445 5355 51503 5361
rect 51445 5352 51457 5355
rect 50856 5324 51457 5352
rect 50856 5312 50862 5324
rect 51445 5321 51457 5324
rect 51491 5321 51503 5355
rect 51445 5315 51503 5321
rect 53193 5355 53251 5361
rect 53193 5321 53205 5355
rect 53239 5352 53251 5355
rect 54110 5352 54116 5364
rect 53239 5324 54116 5352
rect 53239 5321 53251 5324
rect 53193 5315 53251 5321
rect 54110 5312 54116 5324
rect 54168 5312 54174 5364
rect 54846 5312 54852 5364
rect 54904 5352 54910 5364
rect 55306 5352 55312 5364
rect 54904 5324 55312 5352
rect 54904 5312 54910 5324
rect 55306 5312 55312 5324
rect 55364 5352 55370 5364
rect 55953 5355 56011 5361
rect 55953 5352 55965 5355
rect 55364 5324 55965 5352
rect 55364 5312 55370 5324
rect 55953 5321 55965 5324
rect 55999 5321 56011 5355
rect 55953 5315 56011 5321
rect 43714 5244 43720 5296
rect 43772 5244 43778 5296
rect 45554 5244 45560 5296
rect 45612 5284 45618 5296
rect 47854 5284 47860 5296
rect 45612 5256 47164 5284
rect 47815 5256 47860 5284
rect 45612 5244 45618 5256
rect 41555 5188 43116 5216
rect 41555 5185 41567 5188
rect 41509 5179 41567 5185
rect 44634 5176 44640 5228
rect 44692 5216 44698 5228
rect 45278 5216 45284 5228
rect 44692 5188 45284 5216
rect 44692 5176 44698 5188
rect 45278 5176 45284 5188
rect 45336 5176 45342 5228
rect 47026 5216 47032 5228
rect 46987 5188 47032 5216
rect 47026 5176 47032 5188
rect 47084 5176 47090 5228
rect 47136 5216 47164 5256
rect 47854 5244 47860 5256
rect 47912 5244 47918 5296
rect 50522 5284 50528 5296
rect 48516 5256 50528 5284
rect 48516 5216 48544 5256
rect 50522 5244 50528 5256
rect 50580 5244 50586 5296
rect 53742 5244 53748 5296
rect 53800 5284 53806 5296
rect 53837 5287 53895 5293
rect 53837 5284 53849 5287
rect 53800 5256 53849 5284
rect 53800 5244 53806 5256
rect 53837 5253 53849 5256
rect 53883 5253 53895 5287
rect 53837 5247 53895 5253
rect 54941 5287 54999 5293
rect 54941 5253 54953 5287
rect 54987 5284 54999 5287
rect 55122 5284 55128 5296
rect 54987 5256 55128 5284
rect 54987 5253 54999 5256
rect 54941 5247 54999 5253
rect 55122 5244 55128 5256
rect 55180 5244 55186 5296
rect 55493 5287 55551 5293
rect 55493 5253 55505 5287
rect 55539 5284 55551 5287
rect 57974 5284 57980 5296
rect 55539 5256 57980 5284
rect 55539 5253 55551 5256
rect 55493 5247 55551 5253
rect 57974 5244 57980 5256
rect 58032 5244 58038 5296
rect 47136 5188 48544 5216
rect 48590 5176 48596 5228
rect 48648 5216 48654 5228
rect 48869 5219 48927 5225
rect 48869 5216 48881 5219
rect 48648 5188 48881 5216
rect 48648 5176 48654 5188
rect 48869 5185 48881 5188
rect 48915 5216 48927 5219
rect 49326 5216 49332 5228
rect 48915 5188 49188 5216
rect 49287 5188 49332 5216
rect 48915 5185 48927 5188
rect 48869 5179 48927 5185
rect 38010 5148 38016 5160
rect 37844 5120 38016 5148
rect 38010 5108 38016 5120
rect 38068 5108 38074 5160
rect 38562 5148 38568 5160
rect 38523 5120 38568 5148
rect 38562 5108 38568 5120
rect 38620 5108 38626 5160
rect 40586 5148 40592 5160
rect 40547 5120 40592 5148
rect 40586 5108 40592 5120
rect 40644 5108 40650 5160
rect 40954 5108 40960 5160
rect 41012 5148 41018 5160
rect 41598 5148 41604 5160
rect 41012 5120 41604 5148
rect 41012 5108 41018 5120
rect 41598 5108 41604 5120
rect 41656 5108 41662 5160
rect 41693 5151 41751 5157
rect 41693 5117 41705 5151
rect 41739 5148 41751 5151
rect 42058 5148 42064 5160
rect 41739 5120 42064 5148
rect 41739 5117 41751 5120
rect 41693 5111 41751 5117
rect 42058 5108 42064 5120
rect 42116 5108 42122 5160
rect 44361 5151 44419 5157
rect 44361 5148 44373 5151
rect 42904 5120 44373 5148
rect 38930 5080 38936 5092
rect 37292 5052 38936 5080
rect 38930 5040 38936 5052
rect 38988 5040 38994 5092
rect 40770 5040 40776 5092
rect 40828 5080 40834 5092
rect 42904 5080 42932 5120
rect 44361 5117 44373 5120
rect 44407 5117 44419 5151
rect 44361 5111 44419 5117
rect 45830 5108 45836 5160
rect 45888 5148 45894 5160
rect 49050 5148 49056 5160
rect 45888 5120 49056 5148
rect 45888 5108 45894 5120
rect 49050 5108 49056 5120
rect 49108 5108 49114 5160
rect 40828 5052 42932 5080
rect 40828 5040 40834 5052
rect 48498 5040 48504 5092
rect 48556 5080 48562 5092
rect 49160 5080 49188 5188
rect 49326 5176 49332 5188
rect 49384 5176 49390 5228
rect 51626 5216 51632 5228
rect 51587 5188 51632 5216
rect 51626 5176 51632 5188
rect 51684 5176 51690 5228
rect 52270 5176 52276 5228
rect 52328 5216 52334 5228
rect 52365 5219 52423 5225
rect 52365 5216 52377 5219
rect 52328 5188 52377 5216
rect 52328 5176 52334 5188
rect 52365 5185 52377 5188
rect 52411 5185 52423 5219
rect 52365 5179 52423 5185
rect 53285 5219 53343 5225
rect 53285 5185 53297 5219
rect 53331 5216 53343 5219
rect 53466 5216 53472 5228
rect 53331 5188 53472 5216
rect 53331 5185 53343 5188
rect 53285 5179 53343 5185
rect 53466 5176 53472 5188
rect 53524 5176 53530 5228
rect 49234 5108 49240 5160
rect 49292 5148 49298 5160
rect 49513 5151 49571 5157
rect 49513 5148 49525 5151
rect 49292 5120 49525 5148
rect 49292 5108 49298 5120
rect 49513 5117 49525 5120
rect 49559 5117 49571 5151
rect 49513 5111 49571 5117
rect 49602 5108 49608 5160
rect 49660 5148 49666 5160
rect 53760 5148 53788 5244
rect 54573 5219 54631 5225
rect 54573 5185 54585 5219
rect 54619 5185 54631 5219
rect 55140 5216 55168 5244
rect 56042 5216 56048 5228
rect 55140 5188 56048 5216
rect 54573 5179 54631 5185
rect 54588 5148 54616 5179
rect 56042 5176 56048 5188
rect 56100 5216 56106 5228
rect 57057 5219 57115 5225
rect 57057 5216 57069 5219
rect 56100 5188 57069 5216
rect 56100 5176 56106 5188
rect 57057 5185 57069 5188
rect 57103 5185 57115 5219
rect 57057 5179 57115 5185
rect 54662 5148 54668 5160
rect 49660 5120 53788 5148
rect 54575 5120 54668 5148
rect 49660 5108 49666 5120
rect 54662 5108 54668 5120
rect 54720 5148 54726 5160
rect 57514 5148 57520 5160
rect 54720 5120 57520 5148
rect 54720 5108 54726 5120
rect 57514 5108 57520 5120
rect 57572 5108 57578 5160
rect 50614 5080 50620 5092
rect 48556 5052 48912 5080
rect 49160 5052 50620 5080
rect 48556 5040 48562 5052
rect 32364 4984 33272 5012
rect 32364 4972 32370 4984
rect 37274 4972 37280 5024
rect 37332 5012 37338 5024
rect 37553 5015 37611 5021
rect 37553 5012 37565 5015
rect 37332 4984 37565 5012
rect 37332 4972 37338 4984
rect 37553 4981 37565 4984
rect 37599 4981 37611 5015
rect 37553 4975 37611 4981
rect 40494 4972 40500 5024
rect 40552 5012 40558 5024
rect 41049 5015 41107 5021
rect 41049 5012 41061 5015
rect 40552 4984 41061 5012
rect 40552 4972 40558 4984
rect 41049 4981 41061 4984
rect 41095 4981 41107 5015
rect 41049 4975 41107 4981
rect 41598 4972 41604 5024
rect 41656 5012 41662 5024
rect 45097 5015 45155 5021
rect 45097 5012 45109 5015
rect 41656 4984 45109 5012
rect 41656 4972 41662 4984
rect 45097 4981 45109 4984
rect 45143 5012 45155 5015
rect 46198 5012 46204 5024
rect 45143 4984 46204 5012
rect 45143 4981 45155 4984
rect 45097 4975 45155 4981
rect 46198 4972 46204 4984
rect 46256 4972 46262 5024
rect 46293 5015 46351 5021
rect 46293 4981 46305 5015
rect 46339 5012 46351 5015
rect 46474 5012 46480 5024
rect 46339 4984 46480 5012
rect 46339 4981 46351 4984
rect 46293 4975 46351 4981
rect 46474 4972 46480 4984
rect 46532 5012 46538 5024
rect 48590 5012 48596 5024
rect 46532 4984 48596 5012
rect 46532 4972 46538 4984
rect 48590 4972 48596 4984
rect 48648 4972 48654 5024
rect 48774 5012 48780 5024
rect 48735 4984 48780 5012
rect 48774 4972 48780 4984
rect 48832 4972 48838 5024
rect 48884 5012 48912 5052
rect 50614 5040 50620 5052
rect 50672 5080 50678 5092
rect 52181 5083 52239 5089
rect 52181 5080 52193 5083
rect 50672 5052 52193 5080
rect 50672 5040 50678 5052
rect 52181 5049 52193 5052
rect 52227 5049 52239 5083
rect 52181 5043 52239 5049
rect 50798 5012 50804 5024
rect 48884 4984 50804 5012
rect 50798 4972 50804 4984
rect 50856 4972 50862 5024
rect 51626 4972 51632 5024
rect 51684 5012 51690 5024
rect 55030 5012 55036 5024
rect 51684 4984 55036 5012
rect 51684 4972 51690 4984
rect 55030 4972 55036 4984
rect 55088 4972 55094 5024
rect 56502 5012 56508 5024
rect 56463 4984 56508 5012
rect 56502 4972 56508 4984
rect 56560 4972 56566 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 26050 4768 26056 4820
rect 26108 4808 26114 4820
rect 26237 4811 26295 4817
rect 26237 4808 26249 4811
rect 26108 4780 26249 4808
rect 26108 4768 26114 4780
rect 26237 4777 26249 4780
rect 26283 4808 26295 4811
rect 26697 4811 26755 4817
rect 26697 4808 26709 4811
rect 26283 4780 26709 4808
rect 26283 4777 26295 4780
rect 26237 4771 26295 4777
rect 26697 4777 26709 4780
rect 26743 4777 26755 4811
rect 27246 4808 27252 4820
rect 27207 4780 27252 4808
rect 26697 4771 26755 4777
rect 27246 4768 27252 4780
rect 27304 4768 27310 4820
rect 27706 4768 27712 4820
rect 27764 4808 27770 4820
rect 27801 4811 27859 4817
rect 27801 4808 27813 4811
rect 27764 4780 27813 4808
rect 27764 4768 27770 4780
rect 27801 4777 27813 4780
rect 27847 4777 27859 4811
rect 27801 4771 27859 4777
rect 29089 4811 29147 4817
rect 29089 4777 29101 4811
rect 29135 4808 29147 4811
rect 29362 4808 29368 4820
rect 29135 4780 29368 4808
rect 29135 4777 29147 4780
rect 29089 4771 29147 4777
rect 29362 4768 29368 4780
rect 29420 4768 29426 4820
rect 30006 4768 30012 4820
rect 30064 4808 30070 4820
rect 30101 4811 30159 4817
rect 30101 4808 30113 4811
rect 30064 4780 30113 4808
rect 30064 4768 30070 4780
rect 30101 4777 30113 4780
rect 30147 4777 30159 4811
rect 30101 4771 30159 4777
rect 31021 4811 31079 4817
rect 31021 4777 31033 4811
rect 31067 4808 31079 4811
rect 31110 4808 31116 4820
rect 31067 4780 31116 4808
rect 31067 4777 31079 4780
rect 31021 4771 31079 4777
rect 31110 4768 31116 4780
rect 31168 4768 31174 4820
rect 32490 4808 32496 4820
rect 32451 4780 32496 4808
rect 32490 4768 32496 4780
rect 32548 4768 32554 4820
rect 33042 4768 33048 4820
rect 33100 4808 33106 4820
rect 33686 4808 33692 4820
rect 33100 4780 33692 4808
rect 33100 4768 33106 4780
rect 33686 4768 33692 4780
rect 33744 4808 33750 4820
rect 33965 4811 34023 4817
rect 33965 4808 33977 4811
rect 33744 4780 33977 4808
rect 33744 4768 33750 4780
rect 33965 4777 33977 4780
rect 34011 4808 34023 4811
rect 34146 4808 34152 4820
rect 34011 4780 34152 4808
rect 34011 4777 34023 4780
rect 33965 4771 34023 4777
rect 34146 4768 34152 4780
rect 34204 4808 34210 4820
rect 37550 4808 37556 4820
rect 34204 4780 37556 4808
rect 34204 4768 34210 4780
rect 37550 4768 37556 4780
rect 37608 4768 37614 4820
rect 37826 4768 37832 4820
rect 37884 4808 37890 4820
rect 38289 4811 38347 4817
rect 38289 4808 38301 4811
rect 37884 4780 38301 4808
rect 37884 4768 37890 4780
rect 38289 4777 38301 4780
rect 38335 4777 38347 4811
rect 38289 4771 38347 4777
rect 39117 4811 39175 4817
rect 39117 4777 39129 4811
rect 39163 4808 39175 4811
rect 41322 4808 41328 4820
rect 39163 4780 41328 4808
rect 39163 4777 39175 4780
rect 39117 4771 39175 4777
rect 41322 4768 41328 4780
rect 41380 4768 41386 4820
rect 41874 4768 41880 4820
rect 41932 4808 41938 4820
rect 42426 4808 42432 4820
rect 41932 4780 42432 4808
rect 41932 4768 41938 4780
rect 42426 4768 42432 4780
rect 42484 4768 42490 4820
rect 45738 4808 45744 4820
rect 42536 4780 45744 4808
rect 42536 4752 42564 4780
rect 45738 4768 45744 4780
rect 45796 4768 45802 4820
rect 45830 4768 45836 4820
rect 45888 4808 45894 4820
rect 45888 4780 45933 4808
rect 45888 4768 45894 4780
rect 47394 4768 47400 4820
rect 47452 4808 47458 4820
rect 47452 4780 47497 4808
rect 47452 4768 47458 4780
rect 47670 4768 47676 4820
rect 47728 4808 47734 4820
rect 50341 4811 50399 4817
rect 50341 4808 50353 4811
rect 47728 4780 50353 4808
rect 47728 4768 47734 4780
rect 50341 4777 50353 4780
rect 50387 4777 50399 4811
rect 51534 4808 51540 4820
rect 51495 4780 51540 4808
rect 50341 4771 50399 4777
rect 51534 4768 51540 4780
rect 51592 4768 51598 4820
rect 52733 4811 52791 4817
rect 52733 4777 52745 4811
rect 52779 4808 52791 4811
rect 52822 4808 52828 4820
rect 52779 4780 52828 4808
rect 52779 4777 52791 4780
rect 52733 4771 52791 4777
rect 52822 4768 52828 4780
rect 52880 4768 52886 4820
rect 54018 4768 54024 4820
rect 54076 4808 54082 4820
rect 54205 4811 54263 4817
rect 54205 4808 54217 4811
rect 54076 4780 54217 4808
rect 54076 4768 54082 4780
rect 54205 4777 54217 4780
rect 54251 4777 54263 4811
rect 56042 4808 56048 4820
rect 56003 4780 56048 4808
rect 54205 4771 54263 4777
rect 56042 4768 56048 4780
rect 56100 4808 56106 4820
rect 56597 4811 56655 4817
rect 56597 4808 56609 4811
rect 56100 4780 56609 4808
rect 56100 4768 56106 4780
rect 56597 4777 56609 4780
rect 56643 4777 56655 4811
rect 56597 4771 56655 4777
rect 26326 4700 26332 4752
rect 26384 4740 26390 4752
rect 28077 4743 28135 4749
rect 28077 4740 28089 4743
rect 26384 4712 28089 4740
rect 26384 4700 26390 4712
rect 27816 4684 27844 4712
rect 28077 4709 28089 4712
rect 28123 4709 28135 4743
rect 28077 4703 28135 4709
rect 28810 4700 28816 4752
rect 28868 4740 28874 4752
rect 29733 4743 29791 4749
rect 29733 4740 29745 4743
rect 28868 4712 29745 4740
rect 28868 4700 28874 4712
rect 29733 4709 29745 4712
rect 29779 4709 29791 4743
rect 31202 4740 31208 4752
rect 29733 4703 29791 4709
rect 30024 4712 31208 4740
rect 27798 4632 27804 4684
rect 27856 4632 27862 4684
rect 28169 4675 28227 4681
rect 28169 4641 28181 4675
rect 28215 4672 28227 4675
rect 28350 4672 28356 4684
rect 28215 4644 28356 4672
rect 28215 4641 28227 4644
rect 28169 4635 28227 4641
rect 28350 4632 28356 4644
rect 28408 4672 28414 4684
rect 30024 4672 30052 4712
rect 31202 4700 31208 4712
rect 31260 4700 31266 4752
rect 31846 4740 31852 4752
rect 31759 4712 31852 4740
rect 31846 4700 31852 4712
rect 31904 4740 31910 4752
rect 34333 4743 34391 4749
rect 31904 4712 32996 4740
rect 31904 4700 31910 4712
rect 30190 4672 30196 4684
rect 28408 4644 30052 4672
rect 30151 4644 30196 4672
rect 28408 4632 28414 4644
rect 30190 4632 30196 4644
rect 30248 4632 30254 4684
rect 32968 4672 32996 4712
rect 34333 4709 34345 4743
rect 34379 4740 34391 4743
rect 34606 4740 34612 4752
rect 34379 4712 34612 4740
rect 34379 4709 34391 4712
rect 34333 4703 34391 4709
rect 34606 4700 34612 4712
rect 34664 4700 34670 4752
rect 38562 4700 38568 4752
rect 38620 4740 38626 4752
rect 42518 4740 42524 4752
rect 38620 4712 42524 4740
rect 38620 4700 38626 4712
rect 42518 4700 42524 4712
rect 42576 4700 42582 4752
rect 43622 4700 43628 4752
rect 43680 4740 43686 4752
rect 43717 4743 43775 4749
rect 43717 4740 43729 4743
rect 43680 4712 43729 4740
rect 43680 4700 43686 4712
rect 43717 4709 43729 4712
rect 43763 4740 43775 4743
rect 47762 4740 47768 4752
rect 43763 4712 47768 4740
rect 43763 4709 43775 4712
rect 43717 4703 43775 4709
rect 47762 4700 47768 4712
rect 47820 4700 47826 4752
rect 49145 4743 49203 4749
rect 49145 4709 49157 4743
rect 49191 4740 49203 4743
rect 49970 4740 49976 4752
rect 49191 4712 49976 4740
rect 49191 4709 49203 4712
rect 49145 4703 49203 4709
rect 33410 4672 33416 4684
rect 32968 4644 33416 4672
rect 33410 4632 33416 4644
rect 33468 4672 33474 4684
rect 33778 4672 33784 4684
rect 33468 4644 33784 4672
rect 33468 4632 33474 4644
rect 33778 4632 33784 4644
rect 33836 4632 33842 4684
rect 33870 4632 33876 4684
rect 33928 4672 33934 4684
rect 37090 4672 37096 4684
rect 33928 4644 37096 4672
rect 33928 4632 33934 4644
rect 37090 4632 37096 4644
rect 37148 4632 37154 4684
rect 37458 4632 37464 4684
rect 37516 4672 37522 4684
rect 37829 4675 37887 4681
rect 37829 4672 37841 4675
rect 37516 4644 37841 4672
rect 37516 4632 37522 4644
rect 37829 4641 37841 4644
rect 37875 4641 37887 4675
rect 40218 4672 40224 4684
rect 37829 4635 37887 4641
rect 39040 4644 40224 4672
rect 27985 4607 28043 4613
rect 27985 4573 27997 4607
rect 28031 4604 28043 4607
rect 28074 4604 28080 4616
rect 28031 4576 28080 4604
rect 28031 4573 28043 4576
rect 27985 4567 28043 4573
rect 28074 4564 28080 4576
rect 28132 4564 28138 4616
rect 28258 4604 28264 4616
rect 28219 4576 28264 4604
rect 28258 4564 28264 4576
rect 28316 4564 28322 4616
rect 28442 4604 28448 4616
rect 28403 4576 28448 4604
rect 28442 4564 28448 4576
rect 28500 4564 28506 4616
rect 28997 4607 29055 4613
rect 28997 4604 29009 4607
rect 28552 4576 29009 4604
rect 25314 4496 25320 4548
rect 25372 4536 25378 4548
rect 28552 4536 28580 4576
rect 28997 4573 29009 4576
rect 29043 4573 29055 4607
rect 28997 4567 29055 4573
rect 25372 4508 28580 4536
rect 29012 4536 29040 4567
rect 29086 4564 29092 4616
rect 29144 4604 29150 4616
rect 29181 4607 29239 4613
rect 29181 4604 29193 4607
rect 29144 4576 29193 4604
rect 29144 4564 29150 4576
rect 29181 4573 29193 4576
rect 29227 4573 29239 4607
rect 29181 4567 29239 4573
rect 29822 4564 29828 4616
rect 29880 4604 29886 4616
rect 29917 4607 29975 4613
rect 29917 4604 29929 4607
rect 29880 4576 29929 4604
rect 29880 4564 29886 4576
rect 29917 4573 29929 4576
rect 29963 4573 29975 4607
rect 31478 4604 31484 4616
rect 29917 4567 29975 4573
rect 30760 4576 31484 4604
rect 30760 4536 30788 4576
rect 31478 4564 31484 4576
rect 31536 4564 31542 4616
rect 32306 4564 32312 4616
rect 32364 4604 32370 4616
rect 32401 4607 32459 4613
rect 32401 4604 32413 4607
rect 32364 4576 32413 4604
rect 32364 4564 32370 4576
rect 32401 4573 32413 4576
rect 32447 4573 32459 4607
rect 32858 4604 32864 4616
rect 32819 4576 32864 4604
rect 32401 4567 32459 4573
rect 32858 4564 32864 4576
rect 32916 4564 32922 4616
rect 38102 4564 38108 4616
rect 38160 4604 38166 4616
rect 39040 4613 39068 4644
rect 40218 4632 40224 4644
rect 40276 4672 40282 4684
rect 41690 4672 41696 4684
rect 40276 4644 41696 4672
rect 40276 4632 40282 4644
rect 41690 4632 41696 4644
rect 41748 4632 41754 4684
rect 42150 4672 42156 4684
rect 41984 4644 42156 4672
rect 38289 4607 38347 4613
rect 38289 4604 38301 4607
rect 38160 4576 38301 4604
rect 38160 4564 38166 4576
rect 38289 4573 38301 4576
rect 38335 4573 38347 4607
rect 38289 4567 38347 4573
rect 39025 4607 39083 4613
rect 39025 4573 39037 4607
rect 39071 4573 39083 4607
rect 39025 4567 39083 4573
rect 39209 4607 39267 4613
rect 39209 4573 39221 4607
rect 39255 4604 39267 4607
rect 41874 4604 41880 4616
rect 39255 4576 41880 4604
rect 39255 4573 39267 4576
rect 39209 4567 39267 4573
rect 41874 4564 41880 4576
rect 41932 4564 41938 4616
rect 41984 4613 42012 4644
rect 42150 4632 42156 4644
rect 42208 4632 42214 4684
rect 42426 4632 42432 4684
rect 42484 4672 42490 4684
rect 45186 4672 45192 4684
rect 42484 4644 45192 4672
rect 42484 4632 42490 4644
rect 45186 4632 45192 4644
rect 45244 4632 45250 4684
rect 45738 4632 45744 4684
rect 45796 4672 45802 4684
rect 48866 4672 48872 4684
rect 45796 4644 48872 4672
rect 45796 4632 45802 4644
rect 48866 4632 48872 4644
rect 48924 4672 48930 4684
rect 49326 4672 49332 4684
rect 48924 4644 49332 4672
rect 48924 4632 48930 4644
rect 49326 4632 49332 4644
rect 49384 4632 49390 4684
rect 41969 4607 42027 4613
rect 41969 4573 41981 4607
rect 42015 4573 42027 4607
rect 41969 4567 42027 4573
rect 42058 4564 42064 4616
rect 42116 4604 42122 4616
rect 42116 4576 42748 4604
rect 42116 4564 42122 4576
rect 29012 4508 30788 4536
rect 30929 4539 30987 4545
rect 25372 4496 25378 4508
rect 30929 4505 30941 4539
rect 30975 4536 30987 4539
rect 31202 4536 31208 4548
rect 30975 4508 31208 4536
rect 30975 4505 30987 4508
rect 30929 4499 30987 4505
rect 31202 4496 31208 4508
rect 31260 4496 31266 4548
rect 34977 4539 35035 4545
rect 34977 4536 34989 4539
rect 31726 4508 32536 4536
rect 28166 4428 28172 4480
rect 28224 4468 28230 4480
rect 31726 4468 31754 4508
rect 28224 4440 31754 4468
rect 32508 4468 32536 4508
rect 32784 4508 34989 4536
rect 32784 4468 32812 4508
rect 34977 4505 34989 4508
rect 35023 4505 35035 4539
rect 35342 4536 35348 4548
rect 35303 4508 35348 4536
rect 34977 4499 35035 4505
rect 32508 4440 32812 4468
rect 33781 4471 33839 4477
rect 28224 4428 28230 4440
rect 33781 4437 33793 4471
rect 33827 4468 33839 4471
rect 33870 4468 33876 4480
rect 33827 4440 33876 4468
rect 33827 4437 33839 4440
rect 33781 4431 33839 4437
rect 33870 4428 33876 4440
rect 33928 4428 33934 4480
rect 33965 4471 34023 4477
rect 33965 4437 33977 4471
rect 34011 4468 34023 4471
rect 34054 4468 34060 4480
rect 34011 4440 34060 4468
rect 34011 4437 34023 4440
rect 33965 4431 34023 4437
rect 34054 4428 34060 4440
rect 34112 4428 34118 4480
rect 34992 4468 35020 4499
rect 35342 4496 35348 4508
rect 35400 4496 35406 4548
rect 35805 4539 35863 4545
rect 35805 4505 35817 4539
rect 35851 4536 35863 4539
rect 36078 4536 36084 4548
rect 35851 4508 36084 4536
rect 35851 4505 35863 4508
rect 35805 4499 35863 4505
rect 36078 4496 36084 4508
rect 36136 4496 36142 4548
rect 37090 4496 37096 4548
rect 37148 4496 37154 4548
rect 37553 4539 37611 4545
rect 37553 4505 37565 4539
rect 37599 4536 37611 4539
rect 42334 4536 42340 4548
rect 37599 4508 42340 4536
rect 37599 4505 37611 4508
rect 37553 4499 37611 4505
rect 42334 4496 42340 4508
rect 42392 4496 42398 4548
rect 42613 4539 42671 4545
rect 42613 4505 42625 4539
rect 42659 4505 42671 4539
rect 42613 4499 42671 4505
rect 37642 4468 37648 4480
rect 34992 4440 37648 4468
rect 37642 4428 37648 4440
rect 37700 4428 37706 4480
rect 40678 4468 40684 4480
rect 40639 4440 40684 4468
rect 40678 4428 40684 4440
rect 40736 4428 40742 4480
rect 41506 4428 41512 4480
rect 41564 4468 41570 4480
rect 42628 4468 42656 4499
rect 41564 4440 42656 4468
rect 42720 4468 42748 4576
rect 42886 4564 42892 4616
rect 42944 4604 42950 4616
rect 46934 4604 46940 4616
rect 42944 4576 46566 4604
rect 46847 4576 46940 4604
rect 42944 4564 42950 4576
rect 43438 4536 43444 4548
rect 43399 4508 43444 4536
rect 43438 4496 43444 4508
rect 43496 4496 43502 4548
rect 43530 4496 43536 4548
rect 43588 4536 43594 4548
rect 44269 4539 44327 4545
rect 44269 4536 44281 4539
rect 43588 4508 44281 4536
rect 43588 4496 43594 4508
rect 44269 4505 44281 4508
rect 44315 4536 44327 4539
rect 45186 4536 45192 4548
rect 44315 4508 45192 4536
rect 44315 4505 44327 4508
rect 44269 4499 44327 4505
rect 45186 4496 45192 4508
rect 45244 4536 45250 4548
rect 46014 4536 46020 4548
rect 45244 4508 46020 4536
rect 45244 4496 45250 4508
rect 46014 4496 46020 4508
rect 46072 4496 46078 4548
rect 44174 4468 44180 4480
rect 42720 4440 44180 4468
rect 41564 4428 41570 4440
rect 44174 4428 44180 4440
rect 44232 4428 44238 4480
rect 45646 4428 45652 4480
rect 45704 4468 45710 4480
rect 45922 4468 45928 4480
rect 45704 4440 45928 4468
rect 45704 4428 45710 4440
rect 45922 4428 45928 4440
rect 45980 4468 45986 4480
rect 46293 4471 46351 4477
rect 46293 4468 46305 4471
rect 45980 4440 46305 4468
rect 45980 4428 45986 4440
rect 46293 4437 46305 4440
rect 46339 4468 46351 4471
rect 46382 4468 46388 4480
rect 46339 4440 46388 4468
rect 46339 4437 46351 4440
rect 46293 4431 46351 4437
rect 46382 4428 46388 4440
rect 46440 4428 46446 4480
rect 46538 4468 46566 4576
rect 46934 4564 46940 4576
rect 46992 4604 46998 4616
rect 49436 4604 49464 4712
rect 49970 4700 49976 4712
rect 50028 4700 50034 4752
rect 53098 4740 53104 4752
rect 51046 4712 53104 4740
rect 50798 4632 50804 4684
rect 50856 4672 50862 4684
rect 50893 4675 50951 4681
rect 50893 4672 50905 4675
rect 50856 4644 50905 4672
rect 50856 4632 50862 4644
rect 50893 4641 50905 4644
rect 50939 4672 50951 4675
rect 51046 4672 51074 4712
rect 53098 4700 53104 4712
rect 53156 4740 53162 4752
rect 53561 4743 53619 4749
rect 53561 4740 53573 4743
rect 53156 4712 53573 4740
rect 53156 4700 53162 4712
rect 53561 4709 53573 4712
rect 53607 4740 53619 4743
rect 55214 4740 55220 4752
rect 53607 4712 55220 4740
rect 53607 4709 53619 4712
rect 53561 4703 53619 4709
rect 55214 4700 55220 4712
rect 55272 4740 55278 4752
rect 55493 4743 55551 4749
rect 55493 4740 55505 4743
rect 55272 4712 55505 4740
rect 55272 4700 55278 4712
rect 55493 4709 55505 4712
rect 55539 4709 55551 4743
rect 55493 4703 55551 4709
rect 50939 4644 51074 4672
rect 50939 4641 50951 4644
rect 50893 4635 50951 4641
rect 54202 4632 54208 4684
rect 54260 4672 54266 4684
rect 54757 4675 54815 4681
rect 54757 4672 54769 4675
rect 54260 4644 54769 4672
rect 54260 4632 54266 4644
rect 54757 4641 54769 4644
rect 54803 4641 54815 4675
rect 54757 4635 54815 4641
rect 46992 4576 49464 4604
rect 46992 4564 46998 4576
rect 50154 4564 50160 4616
rect 50212 4604 50218 4616
rect 50522 4604 50528 4616
rect 50212 4576 50528 4604
rect 50212 4564 50218 4576
rect 50522 4564 50528 4576
rect 50580 4604 50586 4616
rect 50709 4607 50767 4613
rect 50709 4604 50721 4607
rect 50580 4576 50721 4604
rect 50580 4564 50586 4576
rect 50709 4573 50721 4576
rect 50755 4573 50767 4607
rect 50709 4567 50767 4573
rect 53377 4607 53435 4613
rect 53377 4573 53389 4607
rect 53423 4604 53435 4607
rect 54570 4604 54576 4616
rect 53423 4576 54576 4604
rect 53423 4573 53435 4576
rect 53377 4567 53435 4573
rect 54570 4564 54576 4576
rect 54628 4604 54634 4616
rect 55582 4604 55588 4616
rect 54628 4576 55588 4604
rect 54628 4564 54634 4576
rect 55582 4564 55588 4576
rect 55640 4564 55646 4616
rect 46658 4496 46664 4548
rect 46716 4536 46722 4548
rect 47949 4539 48007 4545
rect 47949 4536 47961 4539
rect 46716 4508 47961 4536
rect 46716 4496 46722 4508
rect 47949 4505 47961 4508
rect 47995 4505 48007 4539
rect 47949 4499 48007 4505
rect 48038 4496 48044 4548
rect 48096 4536 48102 4548
rect 50801 4539 50859 4545
rect 50801 4536 50813 4539
rect 48096 4508 50813 4536
rect 48096 4496 48102 4508
rect 50801 4505 50813 4508
rect 50847 4505 50859 4539
rect 50801 4499 50859 4505
rect 51994 4496 52000 4548
rect 52052 4536 52058 4548
rect 52457 4539 52515 4545
rect 52457 4536 52469 4539
rect 52052 4508 52469 4536
rect 52052 4496 52058 4508
rect 52457 4505 52469 4508
rect 52503 4505 52515 4539
rect 52457 4499 52515 4505
rect 47302 4468 47308 4480
rect 46538 4440 47308 4468
rect 47302 4428 47308 4440
rect 47360 4428 47366 4480
rect 47486 4428 47492 4480
rect 47544 4468 47550 4480
rect 48501 4471 48559 4477
rect 48501 4468 48513 4471
rect 47544 4440 48513 4468
rect 47544 4428 47550 4440
rect 48501 4437 48513 4440
rect 48547 4437 48559 4471
rect 48501 4431 48559 4437
rect 48590 4428 48596 4480
rect 48648 4468 48654 4480
rect 49602 4468 49608 4480
rect 48648 4440 49608 4468
rect 48648 4428 48654 4440
rect 49602 4428 49608 4440
rect 49660 4428 49666 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 28442 4224 28448 4276
rect 28500 4264 28506 4276
rect 31846 4264 31852 4276
rect 28500 4236 31852 4264
rect 28500 4224 28506 4236
rect 31846 4224 31852 4236
rect 31904 4224 31910 4276
rect 32766 4224 32772 4276
rect 32824 4264 32830 4276
rect 33321 4267 33379 4273
rect 33321 4264 33333 4267
rect 32824 4236 33333 4264
rect 32824 4224 32830 4236
rect 33321 4233 33333 4236
rect 33367 4264 33379 4267
rect 33870 4264 33876 4276
rect 33367 4236 33876 4264
rect 33367 4233 33379 4236
rect 33321 4227 33379 4233
rect 33870 4224 33876 4236
rect 33928 4224 33934 4276
rect 34054 4264 34060 4276
rect 34015 4236 34060 4264
rect 34054 4224 34060 4236
rect 34112 4224 34118 4276
rect 34146 4224 34152 4276
rect 34204 4264 34210 4276
rect 34204 4236 34249 4264
rect 34204 4224 34210 4236
rect 34790 4224 34796 4276
rect 34848 4264 34854 4276
rect 35802 4264 35808 4276
rect 34848 4236 35808 4264
rect 34848 4224 34854 4236
rect 35802 4224 35808 4236
rect 35860 4264 35866 4276
rect 37090 4264 37096 4276
rect 35860 4236 37096 4264
rect 35860 4224 35866 4236
rect 29086 4196 29092 4208
rect 29047 4168 29092 4196
rect 29086 4156 29092 4168
rect 29144 4156 29150 4208
rect 29822 4156 29828 4208
rect 29880 4196 29886 4208
rect 31297 4199 31355 4205
rect 31297 4196 31309 4199
rect 29880 4168 31309 4196
rect 29880 4156 29886 4168
rect 31297 4165 31309 4168
rect 31343 4165 31355 4199
rect 32398 4196 32404 4208
rect 32359 4168 32404 4196
rect 31297 4159 31355 4165
rect 32398 4156 32404 4168
rect 32456 4156 32462 4208
rect 34072 4196 34100 4224
rect 32508 4168 34100 4196
rect 34241 4199 34299 4205
rect 32508 4140 32536 4168
rect 34241 4165 34253 4199
rect 34287 4196 34299 4199
rect 34698 4196 34704 4208
rect 34287 4168 34704 4196
rect 34287 4165 34299 4168
rect 34241 4159 34299 4165
rect 28074 4088 28080 4140
rect 28132 4128 28138 4140
rect 28169 4131 28227 4137
rect 28169 4128 28181 4131
rect 28132 4100 28181 4128
rect 28132 4088 28138 4100
rect 28169 4097 28181 4100
rect 28215 4097 28227 4131
rect 28350 4128 28356 4140
rect 28311 4100 28356 4128
rect 28169 4091 28227 4097
rect 28350 4088 28356 4100
rect 28408 4088 28414 4140
rect 28445 4131 28503 4137
rect 28445 4097 28457 4131
rect 28491 4097 28503 4131
rect 30190 4128 30196 4140
rect 30151 4100 30196 4128
rect 28445 4091 28503 4097
rect 27982 4060 27988 4072
rect 27943 4032 27988 4060
rect 27982 4020 27988 4032
rect 28040 4020 28046 4072
rect 28460 4060 28488 4091
rect 30190 4088 30196 4100
rect 30248 4088 30254 4140
rect 30282 4088 30288 4140
rect 30340 4128 30346 4140
rect 30653 4131 30711 4137
rect 30653 4128 30665 4131
rect 30340 4100 30665 4128
rect 30340 4088 30346 4100
rect 30653 4097 30665 4100
rect 30699 4097 30711 4131
rect 30653 4091 30711 4097
rect 31478 4088 31484 4140
rect 31536 4128 31542 4140
rect 31665 4131 31723 4137
rect 31665 4128 31677 4131
rect 31536 4100 31677 4128
rect 31536 4088 31542 4100
rect 31665 4097 31677 4100
rect 31711 4128 31723 4131
rect 32309 4131 32367 4137
rect 32309 4128 32321 4131
rect 31711 4100 32321 4128
rect 31711 4097 31723 4100
rect 31665 4091 31723 4097
rect 32309 4097 32321 4100
rect 32355 4097 32367 4131
rect 32309 4091 32367 4097
rect 32214 4060 32220 4072
rect 28460 4032 32220 4060
rect 32214 4020 32220 4032
rect 32272 4020 32278 4072
rect 32324 4060 32352 4091
rect 32490 4088 32496 4140
rect 32548 4128 32554 4140
rect 32548 4100 32641 4128
rect 32548 4088 32554 4100
rect 32674 4088 32680 4140
rect 32732 4128 32738 4140
rect 33873 4131 33931 4137
rect 32732 4100 32777 4128
rect 32732 4088 32738 4100
rect 33873 4097 33885 4131
rect 33919 4128 33931 4131
rect 33962 4128 33968 4140
rect 33919 4100 33968 4128
rect 33919 4097 33931 4100
rect 33873 4091 33931 4097
rect 33962 4088 33968 4100
rect 34020 4088 34026 4140
rect 32582 4060 32588 4072
rect 32324 4032 32588 4060
rect 32582 4020 32588 4032
rect 32640 4020 32646 4072
rect 32692 4060 32720 4088
rect 34146 4060 34152 4072
rect 32692 4032 34152 4060
rect 34146 4020 34152 4032
rect 34204 4060 34210 4072
rect 34256 4060 34284 4159
rect 34698 4156 34704 4168
rect 34756 4156 34762 4208
rect 36372 4196 36400 4236
rect 37090 4224 37096 4236
rect 37148 4264 37154 4276
rect 37148 4236 39068 4264
rect 37148 4224 37154 4236
rect 36202 4168 36400 4196
rect 36633 4199 36691 4205
rect 36633 4165 36645 4199
rect 36679 4196 36691 4199
rect 37274 4196 37280 4208
rect 36679 4168 37280 4196
rect 36679 4165 36691 4168
rect 36633 4159 36691 4165
rect 37274 4156 37280 4168
rect 37332 4156 37338 4208
rect 39040 4196 39068 4236
rect 40862 4224 40868 4276
rect 40920 4264 40926 4276
rect 43622 4264 43628 4276
rect 40920 4236 43628 4264
rect 40920 4224 40926 4236
rect 43622 4224 43628 4236
rect 43680 4224 43686 4276
rect 46198 4224 46204 4276
rect 46256 4264 46262 4276
rect 53837 4267 53895 4273
rect 46256 4236 53328 4264
rect 46256 4224 46262 4236
rect 40034 4196 40040 4208
rect 38962 4168 40040 4196
rect 40034 4156 40040 4168
rect 40092 4196 40098 4208
rect 40310 4196 40316 4208
rect 40092 4168 40316 4196
rect 40092 4156 40098 4168
rect 40310 4156 40316 4168
rect 40368 4156 40374 4208
rect 41690 4156 41696 4208
rect 41748 4196 41754 4208
rect 41969 4199 42027 4205
rect 41969 4196 41981 4199
rect 41748 4168 41981 4196
rect 41748 4156 41754 4168
rect 41969 4165 41981 4168
rect 42015 4196 42027 4199
rect 43530 4196 43536 4208
rect 42015 4168 43536 4196
rect 42015 4165 42027 4168
rect 41969 4159 42027 4165
rect 43530 4156 43536 4168
rect 43588 4156 43594 4208
rect 43714 4156 43720 4208
rect 43772 4196 43778 4208
rect 45002 4205 45008 4208
rect 44998 4196 45008 4205
rect 43772 4168 43838 4196
rect 44963 4168 45008 4196
rect 43772 4156 43778 4168
rect 44998 4159 45008 4168
rect 45002 4156 45008 4159
rect 45060 4156 45066 4208
rect 47578 4156 47584 4208
rect 47636 4196 47642 4208
rect 48133 4199 48191 4205
rect 47636 4168 47900 4196
rect 47636 4156 47642 4168
rect 41138 4088 41144 4140
rect 41196 4088 41202 4140
rect 42610 4128 42616 4140
rect 42571 4100 42616 4128
rect 42610 4088 42616 4100
rect 42668 4088 42674 4140
rect 43257 4131 43315 4137
rect 43257 4097 43269 4131
rect 43303 4128 43315 4131
rect 43346 4128 43352 4140
rect 43303 4100 43352 4128
rect 43303 4097 43315 4100
rect 43257 4091 43315 4097
rect 43346 4088 43352 4100
rect 43404 4088 43410 4140
rect 45278 4088 45284 4140
rect 45336 4128 45342 4140
rect 45738 4128 45744 4140
rect 45336 4100 45381 4128
rect 45699 4100 45744 4128
rect 45336 4088 45342 4100
rect 45738 4088 45744 4100
rect 45796 4088 45802 4140
rect 47213 4131 47271 4137
rect 47213 4097 47225 4131
rect 47259 4128 47271 4131
rect 47872 4128 47900 4168
rect 48133 4165 48145 4199
rect 48179 4165 48191 4199
rect 48958 4196 48964 4208
rect 48919 4168 48964 4196
rect 48133 4159 48191 4165
rect 48148 4128 48176 4159
rect 48958 4156 48964 4168
rect 49016 4156 49022 4208
rect 49602 4156 49608 4208
rect 49660 4196 49666 4208
rect 52181 4199 52239 4205
rect 52181 4196 52193 4199
rect 49660 4168 52193 4196
rect 49660 4156 49666 4168
rect 52181 4165 52193 4168
rect 52227 4196 52239 4199
rect 52546 4196 52552 4208
rect 52227 4168 52552 4196
rect 52227 4165 52239 4168
rect 52181 4159 52239 4165
rect 52546 4156 52552 4168
rect 52604 4156 52610 4208
rect 53098 4196 53104 4208
rect 53059 4168 53104 4196
rect 53098 4156 53104 4168
rect 53156 4156 53162 4208
rect 53300 4205 53328 4236
rect 53837 4233 53849 4267
rect 53883 4264 53895 4267
rect 54202 4264 54208 4276
rect 53883 4236 54208 4264
rect 53883 4233 53895 4236
rect 53837 4227 53895 4233
rect 54202 4224 54208 4236
rect 54260 4224 54266 4276
rect 54849 4267 54907 4273
rect 54849 4233 54861 4267
rect 54895 4264 54907 4267
rect 55122 4264 55128 4276
rect 54895 4236 55128 4264
rect 54895 4233 54907 4236
rect 54849 4227 54907 4233
rect 55122 4224 55128 4236
rect 55180 4224 55186 4276
rect 53285 4199 53343 4205
rect 53285 4165 53297 4199
rect 53331 4196 53343 4199
rect 54938 4196 54944 4208
rect 53331 4168 54944 4196
rect 53331 4165 53343 4168
rect 53285 4159 53343 4165
rect 54938 4156 54944 4168
rect 54996 4196 55002 4208
rect 55490 4196 55496 4208
rect 54996 4168 55496 4196
rect 54996 4156 55002 4168
rect 55490 4156 55496 4168
rect 55548 4156 55554 4208
rect 47259 4100 47808 4128
rect 47872 4100 48176 4128
rect 48225 4131 48283 4137
rect 47259 4097 47271 4100
rect 47213 4091 47271 4097
rect 34885 4063 34943 4069
rect 34885 4060 34897 4063
rect 34204 4032 34284 4060
rect 34348 4032 34897 4060
rect 34204 4020 34210 4032
rect 27798 3952 27804 4004
rect 27856 3992 27862 4004
rect 28261 3995 28319 4001
rect 28261 3992 28273 3995
rect 27856 3964 28273 3992
rect 27856 3952 27862 3964
rect 28261 3961 28273 3964
rect 28307 3961 28319 3995
rect 28261 3955 28319 3961
rect 29454 3952 29460 4004
rect 29512 3992 29518 4004
rect 29733 3995 29791 4001
rect 29733 3992 29745 3995
rect 29512 3964 29745 3992
rect 29512 3952 29518 3964
rect 29733 3961 29745 3964
rect 29779 3961 29791 3995
rect 29733 3955 29791 3961
rect 30300 3964 31754 3992
rect 30300 3936 30328 3964
rect 30101 3927 30159 3933
rect 30101 3893 30113 3927
rect 30147 3924 30159 3927
rect 30282 3924 30288 3936
rect 30147 3896 30288 3924
rect 30147 3893 30159 3896
rect 30101 3887 30159 3893
rect 30282 3884 30288 3896
rect 30340 3884 30346 3936
rect 31726 3924 31754 3964
rect 33870 3952 33876 4004
rect 33928 3992 33934 4004
rect 34348 3992 34376 4032
rect 34885 4029 34897 4032
rect 34931 4029 34943 4063
rect 36909 4063 36967 4069
rect 34885 4023 34943 4029
rect 35636 4032 36860 4060
rect 33928 3964 34376 3992
rect 33928 3952 33934 3964
rect 31846 3924 31852 3936
rect 31726 3896 31852 3924
rect 31846 3884 31852 3896
rect 31904 3924 31910 3936
rect 33042 3924 33048 3936
rect 31904 3896 33048 3924
rect 31904 3884 31910 3896
rect 33042 3884 33048 3896
rect 33100 3884 33106 3936
rect 34348 3924 34376 3964
rect 34425 3995 34483 4001
rect 34425 3961 34437 3995
rect 34471 3992 34483 3995
rect 35636 3992 35664 4032
rect 34471 3964 35664 3992
rect 36832 3992 36860 4032
rect 36909 4029 36921 4063
rect 36955 4060 36967 4063
rect 37274 4060 37280 4072
rect 36955 4032 37280 4060
rect 36955 4029 36967 4032
rect 36909 4023 36967 4029
rect 37274 4020 37280 4032
rect 37332 4060 37338 4072
rect 37458 4060 37464 4072
rect 37332 4032 37464 4060
rect 37332 4020 37338 4032
rect 37458 4020 37464 4032
rect 37516 4020 37522 4072
rect 37734 4060 37740 4072
rect 37695 4032 37740 4060
rect 37734 4020 37740 4032
rect 37792 4020 37798 4072
rect 38470 4020 38476 4072
rect 38528 4060 38534 4072
rect 39761 4063 39819 4069
rect 39761 4060 39773 4063
rect 38528 4032 39773 4060
rect 38528 4020 38534 4032
rect 39761 4029 39773 4032
rect 39807 4029 39819 4063
rect 40034 4060 40040 4072
rect 39995 4032 40040 4060
rect 39761 4023 39819 4029
rect 40034 4020 40040 4032
rect 40092 4020 40098 4072
rect 41506 3992 41512 4004
rect 36832 3964 37504 3992
rect 41419 3964 41512 3992
rect 34471 3961 34483 3964
rect 34425 3955 34483 3961
rect 37366 3924 37372 3936
rect 34348 3896 37372 3924
rect 37366 3884 37372 3896
rect 37424 3884 37430 3936
rect 37476 3924 37504 3964
rect 41506 3952 41512 3964
rect 41564 3992 41570 4004
rect 41564 3964 43484 3992
rect 41564 3952 41570 3964
rect 43456 3936 43484 3964
rect 45554 3952 45560 4004
rect 45612 3992 45618 4004
rect 47780 4001 47808 4100
rect 48225 4097 48237 4131
rect 48271 4097 48283 4131
rect 48225 4091 48283 4097
rect 49513 4131 49571 4137
rect 49513 4097 49525 4131
rect 49559 4128 49571 4131
rect 49878 4128 49884 4140
rect 49559 4100 49884 4128
rect 49559 4097 49571 4100
rect 49513 4091 49571 4097
rect 46293 3995 46351 4001
rect 46293 3992 46305 3995
rect 45612 3964 46305 3992
rect 45612 3952 45618 3964
rect 46293 3961 46305 3964
rect 46339 3961 46351 3995
rect 46293 3955 46351 3961
rect 47765 3995 47823 4001
rect 47765 3961 47777 3995
rect 47811 3961 47823 3995
rect 47765 3955 47823 3961
rect 48130 3952 48136 4004
rect 48188 3992 48194 4004
rect 48240 3992 48268 4091
rect 49878 4088 49884 4100
rect 49936 4088 49942 4140
rect 50709 4131 50767 4137
rect 50709 4097 50721 4131
rect 50755 4128 50767 4131
rect 50890 4128 50896 4140
rect 50755 4100 50896 4128
rect 50755 4097 50767 4100
rect 50709 4091 50767 4097
rect 50890 4088 50896 4100
rect 50948 4088 50954 4140
rect 48409 4063 48467 4069
rect 48409 4029 48421 4063
rect 48455 4060 48467 4063
rect 52917 4063 52975 4069
rect 52917 4060 52929 4063
rect 48455 4032 52929 4060
rect 48455 4029 48467 4032
rect 48409 4023 48467 4029
rect 52917 4029 52929 4032
rect 52963 4029 52975 4063
rect 52917 4023 52975 4029
rect 54202 4020 54208 4072
rect 54260 4060 54266 4072
rect 55953 4063 56011 4069
rect 55953 4060 55965 4063
rect 54260 4032 55965 4060
rect 54260 4020 54266 4032
rect 55953 4029 55965 4032
rect 55999 4029 56011 4063
rect 55953 4023 56011 4029
rect 48188 3964 48268 3992
rect 50157 3995 50215 4001
rect 48188 3952 48194 3964
rect 50157 3961 50169 3995
rect 50203 3992 50215 3995
rect 50706 3992 50712 4004
rect 50203 3964 50712 3992
rect 50203 3961 50215 3964
rect 50157 3955 50215 3961
rect 50706 3952 50712 3964
rect 50764 3952 50770 4004
rect 52178 3952 52184 4004
rect 52236 3992 52242 4004
rect 54662 3992 54668 4004
rect 52236 3964 54668 3992
rect 52236 3952 52242 3964
rect 54662 3952 54668 3964
rect 54720 3952 54726 4004
rect 38286 3924 38292 3936
rect 37476 3896 38292 3924
rect 38286 3884 38292 3896
rect 38344 3884 38350 3936
rect 39209 3927 39267 3933
rect 39209 3893 39221 3927
rect 39255 3924 39267 3927
rect 43346 3924 43352 3936
rect 39255 3896 43352 3924
rect 39255 3893 39267 3896
rect 39209 3887 39267 3893
rect 43346 3884 43352 3896
rect 43404 3884 43410 3936
rect 43438 3884 43444 3936
rect 43496 3924 43502 3936
rect 45646 3924 45652 3936
rect 43496 3896 45652 3924
rect 43496 3884 43502 3896
rect 45646 3884 45652 3896
rect 45704 3884 45710 3936
rect 46474 3884 46480 3936
rect 46532 3924 46538 3936
rect 47029 3927 47087 3933
rect 47029 3924 47041 3927
rect 46532 3896 47041 3924
rect 46532 3884 46538 3896
rect 47029 3893 47041 3896
rect 47075 3893 47087 3927
rect 47029 3887 47087 3893
rect 48222 3884 48228 3936
rect 48280 3924 48286 3936
rect 51166 3924 51172 3936
rect 48280 3896 51172 3924
rect 48280 3884 48286 3896
rect 51166 3884 51172 3896
rect 51224 3884 51230 3936
rect 53466 3884 53472 3936
rect 53524 3924 53530 3936
rect 54297 3927 54355 3933
rect 54297 3924 54309 3927
rect 53524 3896 54309 3924
rect 53524 3884 53530 3896
rect 54297 3893 54309 3896
rect 54343 3924 54355 3927
rect 55401 3927 55459 3933
rect 55401 3924 55413 3927
rect 54343 3896 55413 3924
rect 54343 3893 54355 3896
rect 54297 3887 54355 3893
rect 55401 3893 55413 3896
rect 55447 3893 55459 3927
rect 55401 3887 55459 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 28442 3680 28448 3732
rect 28500 3720 28506 3732
rect 28537 3723 28595 3729
rect 28537 3720 28549 3723
rect 28500 3692 28549 3720
rect 28500 3680 28506 3692
rect 28537 3689 28549 3692
rect 28583 3689 28595 3723
rect 29730 3720 29736 3732
rect 29691 3692 29736 3720
rect 28537 3683 28595 3689
rect 29730 3680 29736 3692
rect 29788 3680 29794 3732
rect 30006 3680 30012 3732
rect 30064 3720 30070 3732
rect 30929 3723 30987 3729
rect 30929 3720 30941 3723
rect 30064 3692 30941 3720
rect 30064 3680 30070 3692
rect 30929 3689 30941 3692
rect 30975 3689 30987 3723
rect 31294 3720 31300 3732
rect 31255 3692 31300 3720
rect 30929 3683 30987 3689
rect 29917 3587 29975 3593
rect 29917 3553 29929 3587
rect 29963 3584 29975 3587
rect 30024 3584 30052 3680
rect 30944 3652 30972 3683
rect 31294 3680 31300 3692
rect 31352 3680 31358 3732
rect 31846 3720 31852 3732
rect 31807 3692 31852 3720
rect 31846 3680 31852 3692
rect 31904 3680 31910 3732
rect 32214 3680 32220 3732
rect 32272 3720 32278 3732
rect 33597 3723 33655 3729
rect 33597 3720 33609 3723
rect 32272 3692 33609 3720
rect 32272 3680 32278 3692
rect 33597 3689 33609 3692
rect 33643 3689 33655 3723
rect 33597 3683 33655 3689
rect 33686 3680 33692 3732
rect 33744 3720 33750 3732
rect 33781 3723 33839 3729
rect 33781 3720 33793 3723
rect 33744 3692 33793 3720
rect 33744 3680 33750 3692
rect 33781 3689 33793 3692
rect 33827 3689 33839 3723
rect 33781 3683 33839 3689
rect 37182 3680 37188 3732
rect 37240 3720 37246 3732
rect 38657 3723 38715 3729
rect 37240 3692 37596 3720
rect 37240 3680 37246 3692
rect 32674 3652 32680 3664
rect 30944 3624 32680 3652
rect 32674 3612 32680 3624
rect 32732 3612 32738 3664
rect 32858 3612 32864 3664
rect 32916 3652 32922 3664
rect 34054 3652 34060 3664
rect 32916 3624 34060 3652
rect 32916 3612 32922 3624
rect 34054 3612 34060 3624
rect 34112 3652 34118 3664
rect 34977 3655 35035 3661
rect 34977 3652 34989 3655
rect 34112 3624 34989 3652
rect 34112 3612 34118 3624
rect 34977 3621 34989 3624
rect 35023 3652 35035 3655
rect 36262 3652 36268 3664
rect 35023 3624 36268 3652
rect 35023 3621 35035 3624
rect 34977 3615 35035 3621
rect 36262 3612 36268 3624
rect 36320 3612 36326 3664
rect 37568 3652 37596 3692
rect 38657 3689 38669 3723
rect 38703 3720 38715 3723
rect 40034 3720 40040 3732
rect 38703 3692 40040 3720
rect 38703 3689 38715 3692
rect 38657 3683 38715 3689
rect 40034 3680 40040 3692
rect 40092 3680 40098 3732
rect 43346 3680 43352 3732
rect 43404 3720 43410 3732
rect 47578 3720 47584 3732
rect 43404 3692 47440 3720
rect 47539 3692 47584 3720
rect 43404 3680 43410 3692
rect 40313 3655 40371 3661
rect 40313 3652 40325 3655
rect 37568 3624 40325 3652
rect 40313 3621 40325 3624
rect 40359 3621 40371 3655
rect 40313 3615 40371 3621
rect 44269 3655 44327 3661
rect 44269 3621 44281 3655
rect 44315 3652 44327 3655
rect 45738 3652 45744 3664
rect 44315 3624 45744 3652
rect 44315 3621 44327 3624
rect 44269 3615 44327 3621
rect 45738 3612 45744 3624
rect 45796 3612 45802 3664
rect 29963 3556 30052 3584
rect 29963 3553 29975 3556
rect 29917 3547 29975 3553
rect 30282 3544 30288 3596
rect 30340 3584 30346 3596
rect 30377 3587 30435 3593
rect 30377 3584 30389 3587
rect 30340 3556 30389 3584
rect 30340 3544 30346 3556
rect 30377 3553 30389 3556
rect 30423 3553 30435 3587
rect 33962 3584 33968 3596
rect 30377 3547 30435 3553
rect 32692 3556 33968 3584
rect 30009 3519 30067 3525
rect 30009 3485 30021 3519
rect 30055 3516 30067 3519
rect 30190 3516 30196 3528
rect 30055 3488 30196 3516
rect 30055 3485 30067 3488
rect 30009 3479 30067 3485
rect 30190 3476 30196 3488
rect 30248 3516 30254 3528
rect 30837 3519 30895 3525
rect 30837 3516 30849 3519
rect 30248 3488 30849 3516
rect 30248 3476 30254 3488
rect 30837 3485 30849 3488
rect 30883 3516 30895 3519
rect 32401 3519 32459 3525
rect 32401 3516 32413 3519
rect 30883 3488 32413 3516
rect 30883 3485 30895 3488
rect 30837 3479 30895 3485
rect 32401 3485 32413 3488
rect 32447 3516 32459 3519
rect 32490 3516 32496 3528
rect 32447 3488 32496 3516
rect 32447 3485 32459 3488
rect 32401 3479 32459 3485
rect 32490 3476 32496 3488
rect 32548 3476 32554 3528
rect 32582 3476 32588 3528
rect 32640 3525 32646 3528
rect 32640 3519 32655 3525
rect 32643 3516 32655 3519
rect 32692 3516 32720 3556
rect 33962 3544 33968 3556
rect 34020 3584 34026 3596
rect 34241 3587 34299 3593
rect 34241 3584 34253 3587
rect 34020 3556 34253 3584
rect 34020 3544 34026 3556
rect 34241 3553 34253 3556
rect 34287 3553 34299 3587
rect 34241 3547 34299 3553
rect 34330 3544 34336 3596
rect 34388 3584 34394 3596
rect 34388 3556 35664 3584
rect 34388 3544 34394 3556
rect 33781 3519 33839 3525
rect 32643 3488 32733 3516
rect 32643 3485 32655 3488
rect 32640 3479 32655 3485
rect 33781 3485 33793 3519
rect 33827 3516 33839 3519
rect 33870 3516 33876 3528
rect 33827 3488 33876 3516
rect 33827 3485 33839 3488
rect 33781 3479 33839 3485
rect 32640 3476 32646 3479
rect 33870 3476 33876 3488
rect 33928 3476 33934 3528
rect 34054 3476 34060 3528
rect 34112 3516 34118 3528
rect 34149 3519 34207 3525
rect 34149 3516 34161 3519
rect 34112 3488 34161 3516
rect 34112 3476 34118 3488
rect 34149 3485 34161 3488
rect 34195 3485 34207 3519
rect 34149 3479 34207 3485
rect 35161 3519 35219 3525
rect 35161 3485 35173 3519
rect 35207 3485 35219 3519
rect 35161 3479 35219 3485
rect 32309 3451 32367 3457
rect 32309 3417 32321 3451
rect 32355 3417 32367 3451
rect 32309 3411 32367 3417
rect 32769 3451 32827 3457
rect 32769 3417 32781 3451
rect 32815 3448 32827 3451
rect 33594 3448 33600 3460
rect 32815 3420 33600 3448
rect 32815 3417 32827 3420
rect 32769 3411 32827 3417
rect 31202 3340 31208 3392
rect 31260 3380 31266 3392
rect 32324 3380 32352 3411
rect 33594 3408 33600 3420
rect 33652 3408 33658 3460
rect 34238 3408 34244 3460
rect 34296 3448 34302 3460
rect 35176 3448 35204 3479
rect 35636 3457 35664 3556
rect 37274 3544 37280 3596
rect 37332 3584 37338 3596
rect 37645 3587 37703 3593
rect 37645 3584 37657 3587
rect 37332 3556 37657 3584
rect 37332 3544 37338 3556
rect 37645 3553 37657 3556
rect 37691 3553 37703 3587
rect 37645 3547 37703 3553
rect 40586 3544 40592 3596
rect 40644 3584 40650 3596
rect 40957 3587 41015 3593
rect 40957 3584 40969 3587
rect 40644 3556 40969 3584
rect 40644 3544 40650 3556
rect 40957 3553 40969 3556
rect 41003 3553 41015 3587
rect 41230 3584 41236 3596
rect 41191 3556 41236 3584
rect 40957 3547 41015 3553
rect 41230 3544 41236 3556
rect 41288 3544 41294 3596
rect 42610 3544 42616 3596
rect 42668 3584 42674 3596
rect 42981 3587 43039 3593
rect 42981 3584 42993 3587
rect 42668 3556 42993 3584
rect 42668 3544 42674 3556
rect 42981 3553 42993 3556
rect 43027 3553 43039 3587
rect 42981 3547 43039 3553
rect 45278 3544 45284 3596
rect 45336 3584 45342 3596
rect 45833 3587 45891 3593
rect 45833 3584 45845 3587
rect 45336 3556 45845 3584
rect 45336 3544 45342 3556
rect 45833 3553 45845 3556
rect 45879 3553 45891 3587
rect 45833 3547 45891 3553
rect 46109 3587 46167 3593
rect 46109 3553 46121 3587
rect 46155 3584 46167 3587
rect 46474 3584 46480 3596
rect 46155 3556 46480 3584
rect 46155 3553 46167 3556
rect 46109 3547 46167 3553
rect 46474 3544 46480 3556
rect 46532 3544 46538 3596
rect 38473 3519 38531 3525
rect 38473 3485 38485 3519
rect 38519 3516 38531 3519
rect 40310 3516 40316 3528
rect 38519 3488 40316 3516
rect 38519 3485 38531 3488
rect 38473 3479 38531 3485
rect 40310 3476 40316 3488
rect 40368 3476 40374 3528
rect 40494 3516 40500 3528
rect 40455 3488 40500 3516
rect 40494 3476 40500 3488
rect 40552 3476 40558 3528
rect 43530 3516 43536 3528
rect 43443 3488 43536 3516
rect 43530 3476 43536 3488
rect 43588 3516 43594 3528
rect 43806 3516 43812 3528
rect 43588 3488 43812 3516
rect 43588 3476 43594 3488
rect 43806 3476 43812 3488
rect 43864 3476 43870 3528
rect 34296 3420 35204 3448
rect 34296 3408 34302 3420
rect 34606 3380 34612 3392
rect 31260 3352 34612 3380
rect 31260 3340 31266 3352
rect 34606 3340 34612 3352
rect 34664 3340 34670 3392
rect 35176 3380 35204 3420
rect 35621 3451 35679 3457
rect 35621 3417 35633 3451
rect 35667 3448 35679 3451
rect 35710 3448 35716 3460
rect 35667 3420 35716 3448
rect 35667 3417 35679 3420
rect 35621 3411 35679 3417
rect 35710 3408 35716 3420
rect 35768 3408 35774 3460
rect 37090 3448 37096 3460
rect 36938 3420 37096 3448
rect 37090 3408 37096 3420
rect 37148 3408 37154 3460
rect 37369 3451 37427 3457
rect 37369 3417 37381 3451
rect 37415 3417 37427 3451
rect 37369 3411 37427 3417
rect 36354 3380 36360 3392
rect 35176 3352 36360 3380
rect 36354 3340 36360 3352
rect 36412 3340 36418 3392
rect 37384 3380 37412 3411
rect 37458 3408 37464 3460
rect 37516 3448 37522 3460
rect 39117 3451 39175 3457
rect 39117 3448 39129 3451
rect 37516 3420 39129 3448
rect 37516 3408 37522 3420
rect 39117 3417 39129 3420
rect 39163 3417 39175 3451
rect 43714 3448 43720 3460
rect 42458 3420 43720 3448
rect 39117 3411 39175 3417
rect 43714 3408 43720 3420
rect 43772 3408 43778 3460
rect 46658 3408 46664 3460
rect 46716 3408 46722 3460
rect 47412 3448 47440 3692
rect 47578 3680 47584 3692
rect 47636 3680 47642 3732
rect 49329 3723 49387 3729
rect 49329 3689 49341 3723
rect 49375 3720 49387 3723
rect 50062 3720 50068 3732
rect 49375 3692 50068 3720
rect 49375 3689 49387 3692
rect 49329 3683 49387 3689
rect 50062 3680 50068 3692
rect 50120 3680 50126 3732
rect 53653 3723 53711 3729
rect 53653 3689 53665 3723
rect 53699 3720 53711 3723
rect 54202 3720 54208 3732
rect 53699 3692 54208 3720
rect 53699 3689 53711 3692
rect 53653 3683 53711 3689
rect 54202 3680 54208 3692
rect 54260 3680 54266 3732
rect 54662 3720 54668 3732
rect 54623 3692 54668 3720
rect 54662 3680 54668 3692
rect 54720 3680 54726 3732
rect 55490 3720 55496 3732
rect 55451 3692 55496 3720
rect 55490 3680 55496 3692
rect 55548 3680 55554 3732
rect 47854 3612 47860 3664
rect 47912 3652 47918 3664
rect 48041 3655 48099 3661
rect 48041 3652 48053 3655
rect 47912 3624 48053 3652
rect 47912 3612 47918 3624
rect 48041 3621 48053 3624
rect 48087 3621 48099 3655
rect 49234 3652 49240 3664
rect 49195 3624 49240 3652
rect 48041 3615 48099 3621
rect 49234 3612 49240 3624
rect 49292 3612 49298 3664
rect 51166 3612 51172 3664
rect 51224 3652 51230 3664
rect 54113 3655 54171 3661
rect 54113 3652 54125 3655
rect 51224 3624 54125 3652
rect 51224 3612 51230 3624
rect 54113 3621 54125 3624
rect 54159 3652 54171 3655
rect 56502 3652 56508 3664
rect 54159 3624 56508 3652
rect 54159 3621 54171 3624
rect 54113 3615 54171 3621
rect 56502 3612 56508 3624
rect 56560 3612 56566 3664
rect 48866 3516 48872 3528
rect 48827 3488 48872 3516
rect 48866 3476 48872 3488
rect 48924 3516 48930 3528
rect 50341 3519 50399 3525
rect 50341 3516 50353 3519
rect 48924 3488 50353 3516
rect 48924 3476 48930 3488
rect 50341 3485 50353 3488
rect 50387 3516 50399 3519
rect 51442 3516 51448 3528
rect 50387 3488 51448 3516
rect 50387 3485 50399 3488
rect 50341 3479 50399 3485
rect 51442 3476 51448 3488
rect 51500 3476 51506 3528
rect 52181 3519 52239 3525
rect 52181 3485 52193 3519
rect 52227 3485 52239 3519
rect 52181 3479 52239 3485
rect 51350 3448 51356 3460
rect 47412 3420 51356 3448
rect 51350 3408 51356 3420
rect 51408 3408 51414 3460
rect 51994 3408 52000 3460
rect 52052 3408 52058 3460
rect 40126 3380 40132 3392
rect 37384 3352 40132 3380
rect 40126 3340 40132 3352
rect 40184 3340 40190 3392
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45281 3383 45339 3389
rect 45281 3380 45293 3383
rect 44232 3352 45293 3380
rect 44232 3340 44238 3352
rect 45281 3349 45293 3352
rect 45327 3380 45339 3383
rect 45922 3380 45928 3392
rect 45327 3352 45928 3380
rect 45327 3349 45339 3352
rect 45281 3343 45339 3349
rect 45922 3340 45928 3352
rect 45980 3340 45986 3392
rect 49234 3340 49240 3392
rect 49292 3380 49298 3392
rect 52196 3380 52224 3479
rect 52270 3476 52276 3528
rect 52328 3516 52334 3528
rect 52641 3519 52699 3525
rect 52641 3516 52653 3519
rect 52328 3488 52653 3516
rect 52328 3476 52334 3488
rect 52641 3485 52653 3488
rect 52687 3485 52699 3519
rect 52641 3479 52699 3485
rect 53466 3380 53472 3392
rect 49292 3352 53472 3380
rect 49292 3340 49298 3352
rect 53466 3340 53472 3352
rect 53524 3340 53530 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 26418 3136 26424 3188
rect 26476 3176 26482 3188
rect 31021 3179 31079 3185
rect 31021 3176 31033 3179
rect 26476 3148 31033 3176
rect 26476 3136 26482 3148
rect 31021 3145 31033 3148
rect 31067 3145 31079 3179
rect 34330 3176 34336 3188
rect 31021 3139 31079 3145
rect 33980 3148 34336 3176
rect 30190 3108 30196 3120
rect 30151 3080 30196 3108
rect 30190 3068 30196 3080
rect 30248 3068 30254 3120
rect 30409 3111 30467 3117
rect 30409 3077 30421 3111
rect 30455 3108 30467 3111
rect 31202 3108 31208 3120
rect 30455 3080 31208 3108
rect 30455 3077 30467 3080
rect 30409 3071 30467 3077
rect 31202 3068 31208 3080
rect 31260 3068 31266 3120
rect 31478 3108 31484 3120
rect 31439 3080 31484 3108
rect 31478 3068 31484 3080
rect 31536 3068 31542 3120
rect 32401 3111 32459 3117
rect 32401 3108 32413 3111
rect 31956 3080 32413 3108
rect 29178 3040 29184 3052
rect 29091 3012 29184 3040
rect 29178 3000 29184 3012
rect 29236 3040 29242 3052
rect 31956 3040 31984 3080
rect 32401 3077 32413 3080
rect 32447 3108 32459 3111
rect 32674 3108 32680 3120
rect 32447 3080 32680 3108
rect 32447 3077 32459 3080
rect 32401 3071 32459 3077
rect 32674 3068 32680 3080
rect 32732 3068 32738 3120
rect 32858 3117 32864 3120
rect 32815 3111 32864 3117
rect 32815 3077 32827 3111
rect 32861 3077 32864 3111
rect 32815 3071 32864 3077
rect 32858 3068 32864 3071
rect 32916 3068 32922 3120
rect 29236 3012 31984 3040
rect 29236 3000 29242 3012
rect 32030 3000 32036 3052
rect 32088 3040 32094 3052
rect 33045 3043 33103 3049
rect 33045 3040 33057 3043
rect 32088 3012 33057 3040
rect 32088 3000 32094 3012
rect 33045 3009 33057 3012
rect 33091 3009 33103 3043
rect 33980 3040 34008 3148
rect 34330 3136 34336 3148
rect 34388 3136 34394 3188
rect 34514 3136 34520 3188
rect 34572 3176 34578 3188
rect 37274 3176 37280 3188
rect 34572 3148 37280 3176
rect 34572 3136 34578 3148
rect 34790 3068 34796 3120
rect 34848 3068 34854 3120
rect 35345 3111 35403 3117
rect 35345 3077 35357 3111
rect 35391 3108 35403 3111
rect 35434 3108 35440 3120
rect 35391 3080 35440 3108
rect 35391 3077 35403 3080
rect 35345 3071 35403 3077
rect 35434 3068 35440 3080
rect 35492 3068 35498 3120
rect 35636 3049 35664 3148
rect 37274 3136 37280 3148
rect 37332 3136 37338 3188
rect 37553 3179 37611 3185
rect 37553 3145 37565 3179
rect 37599 3176 37611 3179
rect 37642 3176 37648 3188
rect 37599 3148 37648 3176
rect 37599 3145 37611 3148
rect 37553 3139 37611 3145
rect 37642 3136 37648 3148
rect 37700 3136 37706 3188
rect 40310 3136 40316 3188
rect 40368 3176 40374 3188
rect 41325 3179 41383 3185
rect 41325 3176 41337 3179
rect 40368 3148 41337 3176
rect 40368 3136 40374 3148
rect 41325 3145 41337 3148
rect 41371 3145 41383 3179
rect 41782 3176 41788 3188
rect 41743 3148 41788 3176
rect 41325 3139 41383 3145
rect 41782 3136 41788 3148
rect 41840 3136 41846 3188
rect 43714 3136 43720 3188
rect 43772 3176 43778 3188
rect 47762 3176 47768 3188
rect 43772 3148 46704 3176
rect 47723 3148 47768 3176
rect 43772 3136 43778 3148
rect 35710 3068 35716 3120
rect 35768 3108 35774 3120
rect 39025 3111 39083 3117
rect 35768 3080 36584 3108
rect 35768 3068 35774 3080
rect 33045 3003 33103 3009
rect 33152 3012 34008 3040
rect 35621 3043 35679 3049
rect 27890 2932 27896 2984
rect 27948 2972 27954 2984
rect 33152 2972 33180 3012
rect 35621 3009 35633 3043
rect 35667 3009 35679 3043
rect 35621 3003 35679 3009
rect 36262 3000 36268 3052
rect 36320 3040 36326 3052
rect 36449 3043 36507 3049
rect 36449 3040 36461 3043
rect 36320 3012 36461 3040
rect 36320 3000 36326 3012
rect 36449 3009 36461 3012
rect 36495 3009 36507 3043
rect 36449 3003 36507 3009
rect 27948 2944 33180 2972
rect 27948 2932 27954 2944
rect 30466 2864 30472 2916
rect 30524 2904 30530 2916
rect 30561 2907 30619 2913
rect 30561 2904 30573 2907
rect 30524 2876 30573 2904
rect 30524 2864 30530 2876
rect 30561 2873 30573 2876
rect 30607 2873 30619 2907
rect 31202 2904 31208 2916
rect 31163 2876 31208 2904
rect 30561 2867 30619 2873
rect 31202 2864 31208 2876
rect 31260 2864 31266 2916
rect 33873 2907 33931 2913
rect 33873 2873 33885 2907
rect 33919 2904 33931 2907
rect 34238 2904 34244 2916
rect 33919 2876 34244 2904
rect 33919 2873 33931 2876
rect 33873 2867 33931 2873
rect 34238 2864 34244 2876
rect 34296 2864 34302 2916
rect 36265 2907 36323 2913
rect 36265 2873 36277 2907
rect 36311 2904 36323 2907
rect 36446 2904 36452 2916
rect 36311 2876 36452 2904
rect 36311 2873 36323 2876
rect 36265 2867 36323 2873
rect 36446 2864 36452 2876
rect 36504 2864 36510 2916
rect 36556 2904 36584 3080
rect 39025 3077 39037 3111
rect 39071 3108 39083 3111
rect 39298 3108 39304 3120
rect 39071 3080 39304 3108
rect 39071 3077 39083 3080
rect 39025 3071 39083 3077
rect 39298 3068 39304 3080
rect 39356 3068 39362 3120
rect 40402 3108 40408 3120
rect 40250 3080 40408 3108
rect 40402 3068 40408 3080
rect 40460 3068 40466 3120
rect 40586 3068 40592 3120
rect 40644 3108 40650 3120
rect 42889 3111 42947 3117
rect 40644 3080 42656 3108
rect 40644 3068 40650 3080
rect 37274 3000 37280 3052
rect 37332 3040 37338 3052
rect 38470 3040 38476 3052
rect 37332 3012 38476 3040
rect 37332 3000 37338 3012
rect 38470 3000 38476 3012
rect 38528 3040 38534 3052
rect 38749 3043 38807 3049
rect 38749 3040 38761 3043
rect 38528 3012 38761 3040
rect 38528 3000 38534 3012
rect 38749 3009 38761 3012
rect 38795 3009 38807 3043
rect 38749 3003 38807 3009
rect 40862 3000 40868 3052
rect 40920 3040 40926 3052
rect 41693 3043 41751 3049
rect 41693 3040 41705 3043
rect 40920 3012 41705 3040
rect 40920 3000 40926 3012
rect 41693 3009 41705 3012
rect 41739 3009 41751 3043
rect 41693 3003 41751 3009
rect 37550 2932 37556 2984
rect 37608 2972 37614 2984
rect 38013 2975 38071 2981
rect 38013 2972 38025 2975
rect 37608 2944 38025 2972
rect 37608 2932 37614 2944
rect 38013 2941 38025 2944
rect 38059 2972 38071 2975
rect 38102 2972 38108 2984
rect 38059 2944 38108 2972
rect 38059 2941 38071 2944
rect 38013 2935 38071 2941
rect 38102 2932 38108 2944
rect 38160 2932 38166 2984
rect 40218 2972 40224 2984
rect 38212 2944 40224 2972
rect 38212 2904 38240 2944
rect 40218 2932 40224 2944
rect 40276 2932 40282 2984
rect 40770 2972 40776 2984
rect 40683 2944 40776 2972
rect 40770 2932 40776 2944
rect 40828 2932 40834 2984
rect 40954 2932 40960 2984
rect 41012 2972 41018 2984
rect 42628 2981 42656 3080
rect 42889 3077 42901 3111
rect 42935 3108 42947 3111
rect 42978 3108 42984 3120
rect 42935 3080 42984 3108
rect 42935 3077 42947 3080
rect 42889 3071 42947 3077
rect 42978 3068 42984 3080
rect 43036 3068 43042 3120
rect 44192 3108 44220 3148
rect 46676 3120 46704 3148
rect 47762 3136 47768 3148
rect 47820 3136 47826 3188
rect 48869 3179 48927 3185
rect 48869 3176 48881 3179
rect 48286 3148 48881 3176
rect 45278 3108 45284 3120
rect 44114 3080 44220 3108
rect 45112 3080 45284 3108
rect 45112 3049 45140 3080
rect 45278 3068 45284 3080
rect 45336 3068 45342 3120
rect 45370 3068 45376 3120
rect 45428 3108 45434 3120
rect 46658 3108 46664 3120
rect 45428 3080 45473 3108
rect 46598 3080 46664 3108
rect 45428 3068 45434 3080
rect 46658 3068 46664 3080
rect 46716 3068 46722 3120
rect 46750 3068 46756 3120
rect 46808 3108 46814 3120
rect 48130 3108 48136 3120
rect 46808 3080 48136 3108
rect 46808 3068 46814 3080
rect 48130 3068 48136 3080
rect 48188 3108 48194 3120
rect 48286 3108 48314 3148
rect 48869 3145 48881 3148
rect 48915 3145 48927 3179
rect 48869 3139 48927 3145
rect 49513 3179 49571 3185
rect 49513 3145 49525 3179
rect 49559 3176 49571 3179
rect 50890 3176 50896 3188
rect 49559 3148 50896 3176
rect 49559 3145 49571 3148
rect 49513 3139 49571 3145
rect 48406 3108 48412 3120
rect 48188 3080 48314 3108
rect 48367 3080 48412 3108
rect 48188 3068 48194 3080
rect 48406 3068 48412 3080
rect 48464 3068 48470 3120
rect 48774 3068 48780 3120
rect 48832 3108 48838 3120
rect 49528 3108 49556 3139
rect 50890 3136 50896 3148
rect 50948 3136 50954 3188
rect 51442 3136 51448 3188
rect 51500 3176 51506 3188
rect 51902 3176 51908 3188
rect 51500 3148 51908 3176
rect 51500 3136 51506 3148
rect 51902 3136 51908 3148
rect 51960 3176 51966 3188
rect 51997 3179 52055 3185
rect 51997 3176 52009 3179
rect 51960 3148 52009 3176
rect 51960 3136 51966 3148
rect 51997 3145 52009 3148
rect 52043 3176 52055 3179
rect 52270 3176 52276 3188
rect 52043 3148 52276 3176
rect 52043 3145 52055 3148
rect 51997 3139 52055 3145
rect 52270 3136 52276 3148
rect 52328 3176 52334 3188
rect 52917 3179 52975 3185
rect 52917 3176 52929 3179
rect 52328 3148 52929 3176
rect 52328 3136 52334 3148
rect 52917 3145 52929 3148
rect 52963 3145 52975 3179
rect 53466 3176 53472 3188
rect 53427 3148 53472 3176
rect 52917 3139 52975 3145
rect 53466 3136 53472 3148
rect 53524 3136 53530 3188
rect 54113 3179 54171 3185
rect 54113 3145 54125 3179
rect 54159 3176 54171 3179
rect 54202 3176 54208 3188
rect 54159 3148 54208 3176
rect 54159 3145 54171 3148
rect 54113 3139 54171 3145
rect 54202 3136 54208 3148
rect 54260 3136 54266 3188
rect 54570 3176 54576 3188
rect 54531 3148 54576 3176
rect 54570 3136 54576 3148
rect 54628 3136 54634 3188
rect 55214 3176 55220 3188
rect 55175 3148 55220 3176
rect 55214 3136 55220 3148
rect 55272 3136 55278 3188
rect 58158 3136 58164 3188
rect 58216 3176 58222 3188
rect 58253 3179 58311 3185
rect 58253 3176 58265 3179
rect 58216 3148 58265 3176
rect 58216 3136 58222 3148
rect 58253 3145 58265 3148
rect 58299 3145 58311 3179
rect 58253 3139 58311 3145
rect 50154 3108 50160 3120
rect 48832 3080 49556 3108
rect 50115 3080 50160 3108
rect 48832 3068 48838 3080
rect 50154 3068 50160 3080
rect 50212 3068 50218 3120
rect 50706 3108 50712 3120
rect 50667 3080 50712 3108
rect 50706 3068 50712 3080
rect 50764 3068 50770 3120
rect 45097 3043 45155 3049
rect 45097 3040 45109 3043
rect 44100 3012 45109 3040
rect 41877 2975 41935 2981
rect 41877 2972 41889 2975
rect 41012 2944 41889 2972
rect 41012 2932 41018 2944
rect 41877 2941 41889 2944
rect 41923 2941 41935 2975
rect 41877 2935 41935 2941
rect 42613 2975 42671 2981
rect 42613 2941 42625 2975
rect 42659 2972 42671 2975
rect 43254 2972 43260 2984
rect 42659 2944 43260 2972
rect 42659 2941 42671 2944
rect 42613 2935 42671 2941
rect 43254 2932 43260 2944
rect 43312 2972 43318 2984
rect 44100 2972 44128 3012
rect 45097 3009 45109 3012
rect 45143 3009 45155 3043
rect 47210 3040 47216 3052
rect 45097 3003 45155 3009
rect 46952 3012 47216 3040
rect 43312 2944 44128 2972
rect 44637 2975 44695 2981
rect 43312 2932 43318 2944
rect 44637 2941 44649 2975
rect 44683 2972 44695 2975
rect 46952 2972 46980 3012
rect 47210 3000 47216 3012
rect 47268 3040 47274 3052
rect 48222 3040 48228 3052
rect 47268 3012 48228 3040
rect 47268 3000 47274 3012
rect 48222 3000 48228 3012
rect 48280 3000 48286 3052
rect 51350 3000 51356 3052
rect 51408 3040 51414 3052
rect 51445 3043 51503 3049
rect 51445 3040 51457 3043
rect 51408 3012 51457 3040
rect 51408 3000 51414 3012
rect 51445 3009 51457 3012
rect 51491 3040 51503 3043
rect 52178 3040 52184 3052
rect 51491 3012 52184 3040
rect 51491 3009 51503 3012
rect 51445 3003 51503 3009
rect 52178 3000 52184 3012
rect 52236 3000 52242 3052
rect 47118 2972 47124 2984
rect 44683 2944 46980 2972
rect 47079 2944 47124 2972
rect 44683 2941 44695 2944
rect 44637 2935 44695 2941
rect 47118 2932 47124 2944
rect 47176 2932 47182 2984
rect 36556 2876 38240 2904
rect 29733 2839 29791 2845
rect 29733 2805 29745 2839
rect 29779 2836 29791 2839
rect 30282 2836 30288 2848
rect 29779 2808 30288 2836
rect 29779 2805 29791 2808
rect 29733 2799 29791 2805
rect 30282 2796 30288 2808
rect 30340 2836 30346 2848
rect 30377 2839 30435 2845
rect 30377 2836 30389 2839
rect 30340 2808 30389 2836
rect 30340 2796 30346 2808
rect 30377 2805 30389 2808
rect 30423 2805 30435 2839
rect 30377 2799 30435 2805
rect 31018 2796 31024 2848
rect 31076 2836 31082 2848
rect 32306 2836 32312 2848
rect 31076 2808 32312 2836
rect 31076 2796 31082 2808
rect 32306 2796 32312 2808
rect 32364 2836 32370 2848
rect 32769 2839 32827 2845
rect 32769 2836 32781 2839
rect 32364 2808 32781 2836
rect 32364 2796 32370 2808
rect 32769 2805 32781 2808
rect 32815 2836 32827 2839
rect 33686 2836 33692 2848
rect 32815 2808 33692 2836
rect 32815 2805 32827 2808
rect 32769 2799 32827 2805
rect 33686 2796 33692 2808
rect 33744 2796 33750 2848
rect 36354 2796 36360 2848
rect 36412 2836 36418 2848
rect 40034 2836 40040 2848
rect 36412 2808 40040 2836
rect 36412 2796 36418 2808
rect 40034 2796 40040 2808
rect 40092 2796 40098 2848
rect 40788 2836 40816 2932
rect 42886 2836 42892 2848
rect 40788 2808 42892 2836
rect 42886 2796 42892 2808
rect 42944 2796 42950 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 29178 2632 29184 2644
rect 29139 2604 29184 2632
rect 29178 2592 29184 2604
rect 29236 2592 29242 2644
rect 30193 2635 30251 2641
rect 30193 2601 30205 2635
rect 30239 2632 30251 2635
rect 31018 2632 31024 2644
rect 30239 2604 31024 2632
rect 30239 2601 30251 2604
rect 30193 2595 30251 2601
rect 31018 2592 31024 2604
rect 31076 2592 31082 2644
rect 31113 2635 31171 2641
rect 31113 2601 31125 2635
rect 31159 2632 31171 2635
rect 31159 2604 31248 2632
rect 31159 2601 31171 2604
rect 31113 2595 31171 2601
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 22186 2564 22192 2576
rect 2455 2536 22192 2564
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 2424 2428 2452 2527
rect 22186 2524 22192 2536
rect 22244 2524 22250 2576
rect 30745 2567 30803 2573
rect 30745 2564 30757 2567
rect 29748 2536 30757 2564
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 21358 2496 21364 2508
rect 5767 2468 21364 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 21358 2456 21364 2468
rect 21416 2456 21422 2508
rect 1903 2400 2452 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 5592 2400 6009 2428
rect 5592 2388 5598 2400
rect 5997 2397 6009 2400
rect 6043 2428 6055 2431
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6043 2400 6561 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12434 2428 12440 2440
rect 12023 2400 12440 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2428 17187 2431
rect 22281 2431 22339 2437
rect 17175 2400 17724 2428
rect 17175 2397 17187 2400
rect 17129 2391 17187 2397
rect 17696 2304 17724 2400
rect 22281 2397 22293 2431
rect 22327 2428 22339 2431
rect 28077 2431 28135 2437
rect 22327 2400 22876 2428
rect 22327 2397 22339 2400
rect 22281 2391 22339 2397
rect 22848 2304 22876 2400
rect 28077 2397 28089 2431
rect 28123 2428 28135 2431
rect 28123 2400 28672 2428
rect 28123 2397 28135 2400
rect 28077 2391 28135 2397
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 72 2264 1685 2292
rect 72 2252 78 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11020 2264 11805 2292
rect 11020 2252 11026 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16945 2295 17003 2301
rect 16945 2292 16957 2295
rect 16816 2264 16957 2292
rect 16816 2252 16822 2264
rect 16945 2261 16957 2264
rect 16991 2261 17003 2295
rect 17678 2292 17684 2304
rect 17639 2264 17684 2292
rect 16945 2255 17003 2261
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22097 2295 22155 2301
rect 22097 2292 22109 2295
rect 21968 2264 22109 2292
rect 21968 2252 21974 2264
rect 22097 2261 22109 2264
rect 22143 2261 22155 2295
rect 22830 2292 22836 2304
rect 22791 2264 22836 2292
rect 22097 2255 22155 2261
rect 22830 2252 22836 2264
rect 22888 2252 22894 2304
rect 27706 2252 27712 2304
rect 27764 2292 27770 2304
rect 28644 2301 28672 2400
rect 28902 2388 28908 2440
rect 28960 2428 28966 2440
rect 29748 2428 29776 2536
rect 30745 2533 30757 2536
rect 30791 2533 30803 2567
rect 31220 2564 31248 2604
rect 31294 2592 31300 2644
rect 31352 2632 31358 2644
rect 36262 2632 36268 2644
rect 31352 2604 36268 2632
rect 31352 2592 31358 2604
rect 36262 2592 36268 2604
rect 36320 2592 36326 2644
rect 36817 2635 36875 2641
rect 36817 2601 36829 2635
rect 36863 2632 36875 2635
rect 38102 2632 38108 2644
rect 36863 2604 38108 2632
rect 36863 2601 36875 2604
rect 36817 2595 36875 2601
rect 38102 2592 38108 2604
rect 38160 2632 38166 2644
rect 40865 2635 40923 2641
rect 40865 2632 40877 2635
rect 38160 2604 40877 2632
rect 38160 2592 38166 2604
rect 40865 2601 40877 2604
rect 40911 2632 40923 2635
rect 41322 2632 41328 2644
rect 40911 2604 41328 2632
rect 40911 2601 40923 2604
rect 40865 2595 40923 2601
rect 41322 2592 41328 2604
rect 41380 2592 41386 2644
rect 43162 2592 43168 2644
rect 43220 2632 43226 2644
rect 43901 2635 43959 2641
rect 43901 2632 43913 2635
rect 43220 2604 43913 2632
rect 43220 2592 43226 2604
rect 43901 2601 43913 2604
rect 43947 2601 43959 2635
rect 43901 2595 43959 2601
rect 45186 2592 45192 2644
rect 45244 2632 45250 2644
rect 45281 2635 45339 2641
rect 45281 2632 45293 2635
rect 45244 2604 45293 2632
rect 45244 2592 45250 2604
rect 45281 2601 45293 2604
rect 45327 2601 45339 2635
rect 45281 2595 45339 2601
rect 46198 2592 46204 2644
rect 46256 2632 46262 2644
rect 46385 2635 46443 2641
rect 46385 2632 46397 2635
rect 46256 2604 46397 2632
rect 46256 2592 46262 2604
rect 46385 2601 46397 2604
rect 46431 2601 46443 2635
rect 47026 2632 47032 2644
rect 46987 2604 47032 2632
rect 46385 2595 46443 2601
rect 47026 2592 47032 2604
rect 47084 2592 47090 2644
rect 48409 2635 48467 2641
rect 48409 2601 48421 2635
rect 48455 2632 48467 2635
rect 48682 2632 48688 2644
rect 48455 2604 48688 2632
rect 48455 2601 48467 2604
rect 48409 2595 48467 2601
rect 48682 2592 48688 2604
rect 48740 2592 48746 2644
rect 48866 2632 48872 2644
rect 48827 2604 48872 2632
rect 48866 2592 48872 2604
rect 48924 2592 48930 2644
rect 50890 2592 50896 2644
rect 50948 2632 50954 2644
rect 51077 2635 51135 2641
rect 51077 2632 51089 2635
rect 50948 2604 51089 2632
rect 50948 2592 50954 2604
rect 51077 2601 51089 2604
rect 51123 2601 51135 2635
rect 51626 2632 51632 2644
rect 51587 2604 51632 2632
rect 51077 2595 51135 2601
rect 51626 2592 51632 2604
rect 51684 2592 51690 2644
rect 51902 2592 51908 2644
rect 51960 2632 51966 2644
rect 52181 2635 52239 2641
rect 52181 2632 52193 2635
rect 51960 2604 52193 2632
rect 51960 2592 51966 2604
rect 52181 2601 52193 2604
rect 52227 2632 52239 2635
rect 52917 2635 52975 2641
rect 52917 2632 52929 2635
rect 52227 2604 52929 2632
rect 52227 2601 52239 2604
rect 52181 2595 52239 2601
rect 52917 2601 52929 2604
rect 52963 2601 52975 2635
rect 53466 2632 53472 2644
rect 53427 2604 53472 2632
rect 52917 2595 52975 2601
rect 53466 2592 53472 2604
rect 53524 2592 53530 2644
rect 56962 2632 56968 2644
rect 56923 2604 56968 2632
rect 56962 2592 56968 2604
rect 57020 2592 57026 2644
rect 32401 2567 32459 2573
rect 32401 2564 32413 2567
rect 31220 2536 32413 2564
rect 30745 2527 30803 2533
rect 32401 2533 32413 2536
rect 32447 2564 32459 2567
rect 32490 2564 32496 2576
rect 32447 2536 32496 2564
rect 32447 2533 32459 2536
rect 32401 2527 32459 2533
rect 32490 2524 32496 2536
rect 32548 2524 32554 2576
rect 33870 2524 33876 2576
rect 33928 2564 33934 2576
rect 34057 2567 34115 2573
rect 34057 2564 34069 2567
rect 33928 2536 34069 2564
rect 33928 2524 33934 2536
rect 34057 2533 34069 2536
rect 34103 2533 34115 2567
rect 34057 2527 34115 2533
rect 34790 2524 34796 2576
rect 34848 2564 34854 2576
rect 35161 2567 35219 2573
rect 35161 2564 35173 2567
rect 34848 2536 35173 2564
rect 34848 2524 34854 2536
rect 35161 2533 35173 2536
rect 35207 2533 35219 2567
rect 41877 2567 41935 2573
rect 41877 2564 41889 2567
rect 35161 2527 35219 2533
rect 36280 2536 41889 2564
rect 32508 2496 32536 2524
rect 32508 2468 33640 2496
rect 28960 2400 29776 2428
rect 28960 2388 28966 2400
rect 29914 2388 29920 2440
rect 29972 2428 29978 2440
rect 30009 2431 30067 2437
rect 30009 2428 30021 2431
rect 29972 2400 30021 2428
rect 29972 2388 29978 2400
rect 30009 2397 30021 2400
rect 30055 2397 30067 2431
rect 31202 2428 31208 2440
rect 31163 2400 31208 2428
rect 30009 2391 30067 2397
rect 30024 2360 30052 2391
rect 31202 2388 31208 2400
rect 31260 2388 31266 2440
rect 32585 2431 32643 2437
rect 32585 2397 32597 2431
rect 32631 2428 32643 2431
rect 32674 2428 32680 2440
rect 32631 2400 32680 2428
rect 32631 2397 32643 2400
rect 32585 2391 32643 2397
rect 32674 2388 32680 2400
rect 32732 2388 32738 2440
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33612 2437 33640 2468
rect 33321 2431 33379 2437
rect 33321 2428 33333 2431
rect 33192 2400 33333 2428
rect 33192 2388 33198 2400
rect 33321 2397 33333 2400
rect 33367 2397 33379 2431
rect 33321 2391 33379 2397
rect 33597 2431 33655 2437
rect 33597 2397 33609 2431
rect 33643 2397 33655 2431
rect 34146 2428 34152 2440
rect 34107 2400 34152 2428
rect 33597 2391 33655 2397
rect 34146 2388 34152 2400
rect 34204 2388 34210 2440
rect 35342 2388 35348 2440
rect 35400 2428 35406 2440
rect 36280 2437 36308 2536
rect 41877 2533 41889 2536
rect 41923 2533 41935 2567
rect 43530 2564 43536 2576
rect 41877 2527 41935 2533
rect 42168 2536 43536 2564
rect 37458 2496 37464 2508
rect 37419 2468 37464 2496
rect 37458 2456 37464 2468
rect 37516 2456 37522 2508
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 39132 2468 41429 2496
rect 35437 2431 35495 2437
rect 35437 2428 35449 2431
rect 35400 2400 35449 2428
rect 35400 2388 35406 2400
rect 35437 2397 35449 2400
rect 35483 2428 35495 2431
rect 36265 2431 36323 2437
rect 35483 2400 35894 2428
rect 35483 2397 35495 2400
rect 35437 2391 35495 2397
rect 30024 2332 31800 2360
rect 27893 2295 27951 2301
rect 27893 2292 27905 2295
rect 27764 2264 27905 2292
rect 27764 2252 27770 2264
rect 27893 2261 27905 2264
rect 27939 2261 27951 2295
rect 27893 2255 27951 2261
rect 28629 2295 28687 2301
rect 28629 2261 28641 2295
rect 28675 2292 28687 2295
rect 31294 2292 31300 2304
rect 28675 2264 31300 2292
rect 28675 2261 28687 2264
rect 28629 2255 28687 2261
rect 31294 2252 31300 2264
rect 31352 2252 31358 2304
rect 31772 2301 31800 2332
rect 33502 2320 33508 2372
rect 33560 2360 33566 2372
rect 35866 2360 35894 2400
rect 36265 2397 36277 2431
rect 36311 2397 36323 2431
rect 36265 2391 36323 2397
rect 39132 2360 39160 2468
rect 41417 2465 41429 2468
rect 41463 2496 41475 2499
rect 42168 2496 42196 2536
rect 43530 2524 43536 2536
rect 43588 2524 43594 2576
rect 45646 2524 45652 2576
rect 45704 2564 45710 2576
rect 45833 2567 45891 2573
rect 45833 2564 45845 2567
rect 45704 2536 45845 2564
rect 45704 2524 45710 2536
rect 45833 2533 45845 2536
rect 45879 2533 45891 2567
rect 45833 2527 45891 2533
rect 47118 2524 47124 2576
rect 47176 2564 47182 2576
rect 49234 2564 49240 2576
rect 47176 2536 49240 2564
rect 47176 2524 47182 2536
rect 49234 2524 49240 2536
rect 49292 2564 49298 2576
rect 49421 2567 49479 2573
rect 49421 2564 49433 2567
rect 49292 2536 49433 2564
rect 49292 2524 49298 2536
rect 49421 2533 49433 2536
rect 49467 2533 49479 2567
rect 49421 2527 49479 2533
rect 41463 2468 42196 2496
rect 41463 2465 41475 2468
rect 41417 2459 41475 2465
rect 42242 2456 42248 2508
rect 42300 2496 42306 2508
rect 42300 2468 50660 2496
rect 42300 2456 42306 2468
rect 40034 2428 40040 2440
rect 39995 2400 40040 2428
rect 40034 2388 40040 2400
rect 40092 2388 40098 2440
rect 42061 2431 42119 2437
rect 42061 2397 42073 2431
rect 42107 2428 42119 2431
rect 47026 2428 47032 2440
rect 42107 2400 47032 2428
rect 42107 2397 42119 2400
rect 42061 2391 42119 2397
rect 47026 2388 47032 2400
rect 47084 2388 47090 2440
rect 50632 2437 50660 2468
rect 50617 2431 50675 2437
rect 50617 2397 50629 2431
rect 50663 2428 50675 2431
rect 54021 2431 54079 2437
rect 54021 2428 54033 2431
rect 50663 2400 54033 2428
rect 50663 2397 50675 2400
rect 50617 2391 50675 2397
rect 54021 2397 54033 2400
rect 54067 2397 54079 2431
rect 54021 2391 54079 2397
rect 56413 2431 56471 2437
rect 56413 2397 56425 2431
rect 56459 2428 56471 2431
rect 56962 2428 56968 2440
rect 56459 2400 56968 2428
rect 56459 2397 56471 2400
rect 56413 2391 56471 2397
rect 56962 2388 56968 2400
rect 57020 2388 57026 2440
rect 58069 2431 58127 2437
rect 58069 2397 58081 2431
rect 58115 2428 58127 2431
rect 58158 2428 58164 2440
rect 58115 2400 58164 2428
rect 58115 2397 58127 2400
rect 58069 2391 58127 2397
rect 58158 2388 58164 2400
rect 58216 2388 58222 2440
rect 33560 2332 35296 2360
rect 35866 2332 39160 2360
rect 39209 2363 39267 2369
rect 33560 2320 33566 2332
rect 31757 2295 31815 2301
rect 31757 2261 31769 2295
rect 31803 2292 31815 2295
rect 34422 2292 34428 2304
rect 31803 2264 34428 2292
rect 31803 2261 31815 2264
rect 31757 2255 31815 2261
rect 34422 2252 34428 2264
rect 34480 2252 34486 2304
rect 35268 2292 35296 2332
rect 39209 2329 39221 2363
rect 39255 2360 39267 2363
rect 40678 2360 40684 2372
rect 39255 2332 40684 2360
rect 39255 2329 39267 2332
rect 39209 2323 39267 2329
rect 40678 2320 40684 2332
rect 40736 2360 40742 2372
rect 42613 2363 42671 2369
rect 42613 2360 42625 2363
rect 40736 2332 42625 2360
rect 40736 2320 40742 2332
rect 42613 2329 42625 2332
rect 42659 2329 42671 2363
rect 42613 2323 42671 2329
rect 43530 2320 43536 2372
rect 43588 2360 43594 2372
rect 47765 2363 47823 2369
rect 47765 2360 47777 2363
rect 43588 2332 47777 2360
rect 43588 2320 43594 2332
rect 47765 2329 47777 2332
rect 47811 2329 47823 2363
rect 47765 2323 47823 2329
rect 36081 2295 36139 2301
rect 36081 2292 36093 2295
rect 35268 2264 36093 2292
rect 36081 2261 36093 2264
rect 36127 2261 36139 2295
rect 36081 2255 36139 2261
rect 38654 2252 38660 2304
rect 38712 2292 38718 2304
rect 40221 2295 40279 2301
rect 40221 2292 40233 2295
rect 38712 2264 40233 2292
rect 38712 2252 38718 2264
rect 40221 2261 40233 2264
rect 40267 2261 40279 2295
rect 40221 2255 40279 2261
rect 50154 2252 50160 2304
rect 50212 2292 50218 2304
rect 50433 2295 50491 2301
rect 50433 2292 50445 2295
rect 50212 2264 50445 2292
rect 50212 2252 50218 2264
rect 50433 2261 50445 2264
rect 50479 2261 50491 2295
rect 50433 2255 50491 2261
rect 56042 2252 56048 2304
rect 56100 2292 56106 2304
rect 56229 2295 56287 2301
rect 56229 2292 56241 2295
rect 56100 2264 56241 2292
rect 56100 2252 56106 2264
rect 56229 2261 56241 2264
rect 56275 2261 56287 2295
rect 56229 2255 56287 2261
rect 58253 2295 58311 2301
rect 58253 2261 58265 2295
rect 58299 2292 58311 2295
rect 59906 2292 59912 2304
rect 58299 2264 59912 2292
rect 58299 2261 58311 2264
rect 58253 2255 58311 2261
rect 59906 2252 59912 2264
rect 59964 2252 59970 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 17678 2048 17684 2100
rect 17736 2088 17742 2100
rect 47118 2088 47124 2100
rect 17736 2060 47124 2088
rect 17736 2048 17742 2060
rect 47118 2048 47124 2060
rect 47176 2048 47182 2100
rect 22830 1980 22836 2032
rect 22888 2020 22894 2032
rect 38562 2020 38568 2032
rect 22888 1992 38568 2020
rect 22888 1980 22894 1992
rect 38562 1980 38568 1992
rect 38620 1980 38626 2032
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 2780 57536 2832 57588
rect 3884 57536 3936 57588
rect 9680 57536 9732 57588
rect 15476 57536 15528 57588
rect 21272 57536 21324 57588
rect 26424 57536 26476 57588
rect 38016 57536 38068 57588
rect 43168 57536 43220 57588
rect 48964 57536 49016 57588
rect 54760 57536 54812 57588
rect 58256 57579 58308 57588
rect 58256 57545 58265 57579
rect 58265 57545 58299 57579
rect 58299 57545 58308 57579
rect 58256 57536 58308 57545
rect 28724 57468 28776 57520
rect 2320 57400 2372 57452
rect 4712 57400 4764 57452
rect 10048 57443 10100 57452
rect 10048 57409 10057 57443
rect 10057 57409 10091 57443
rect 10091 57409 10100 57443
rect 10048 57400 10100 57409
rect 15936 57400 15988 57452
rect 22652 57400 22704 57452
rect 27988 57400 28040 57452
rect 32220 57400 32272 57452
rect 43720 57400 43772 57452
rect 49240 57400 49292 57452
rect 55496 57443 55548 57452
rect 55496 57409 55505 57443
rect 55505 57409 55539 57443
rect 55539 57409 55548 57443
rect 55496 57400 55548 57409
rect 57704 57400 57756 57452
rect 32036 57332 32088 57384
rect 2320 57239 2372 57248
rect 2320 57205 2329 57239
rect 2329 57205 2363 57239
rect 2363 57205 2372 57239
rect 2320 57196 2372 57205
rect 4712 57239 4764 57248
rect 4712 57205 4721 57239
rect 4721 57205 4755 57239
rect 4755 57205 4764 57239
rect 4712 57196 4764 57205
rect 22652 57196 22704 57248
rect 27988 57239 28040 57248
rect 27988 57205 27997 57239
rect 27997 57205 28031 57239
rect 28031 57205 28040 57239
rect 27988 57196 28040 57205
rect 43720 57196 43772 57248
rect 57704 57196 57756 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 40408 56788 40460 56840
rect 15936 56695 15988 56704
rect 15936 56661 15945 56695
rect 15945 56661 15979 56695
rect 15979 56661 15988 56695
rect 15936 56652 15988 56661
rect 55496 56720 55548 56772
rect 49240 56652 49292 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 57336 54476 57388 54528
rect 58256 54519 58308 54528
rect 58256 54485 58265 54519
rect 58265 54485 58299 54519
rect 58299 54485 58308 54519
rect 58256 54476 58308 54485
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 1676 53431 1728 53440
rect 1676 53397 1685 53431
rect 1685 53397 1719 53431
rect 1719 53397 1728 53431
rect 1676 53388 1728 53397
rect 2412 53431 2464 53440
rect 2412 53397 2421 53431
rect 2421 53397 2455 53431
rect 2455 53397 2464 53431
rect 2412 53388 2464 53397
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 57796 48696 57848 48748
rect 57796 48492 57848 48544
rect 58256 48535 58308 48544
rect 58256 48501 58265 48535
rect 58265 48501 58299 48535
rect 58299 48501 58308 48535
rect 58256 48492 58308 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 1676 47175 1728 47184
rect 1676 47141 1685 47175
rect 1685 47141 1719 47175
rect 1719 47141 1728 47175
rect 1676 47132 1728 47141
rect 2504 46928 2556 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 57520 42551 57572 42560
rect 57520 42517 57529 42551
rect 57529 42517 57563 42551
rect 57563 42517 57572 42551
rect 57520 42508 57572 42517
rect 58256 42551 58308 42560
rect 58256 42517 58265 42551
rect 58265 42517 58299 42551
rect 58299 42517 58308 42551
rect 58256 42508 58308 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 1860 41123 1912 41132
rect 1860 41089 1869 41123
rect 1869 41089 1903 41123
rect 1903 41089 1912 41123
rect 1860 41080 1912 41089
rect 1676 40919 1728 40928
rect 1676 40885 1685 40919
rect 1685 40885 1719 40919
rect 1719 40885 1728 40919
rect 1676 40876 1728 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 57980 37204 58032 37256
rect 58256 37111 58308 37120
rect 58256 37077 58265 37111
rect 58265 37077 58299 37111
rect 58299 37077 58308 37111
rect 58256 37068 58308 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 1952 35640 2004 35692
rect 1676 35479 1728 35488
rect 1676 35445 1685 35479
rect 1685 35445 1719 35479
rect 1719 35445 1728 35479
rect 1676 35436 1728 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 44824 31331 44876 31340
rect 44824 31297 44833 31331
rect 44833 31297 44867 31331
rect 44867 31297 44876 31331
rect 44824 31288 44876 31297
rect 44916 31288 44968 31340
rect 46756 31331 46808 31340
rect 46756 31297 46765 31331
rect 46765 31297 46799 31331
rect 46799 31297 46808 31331
rect 46756 31288 46808 31297
rect 47032 31331 47084 31340
rect 47032 31297 47041 31331
rect 47041 31297 47075 31331
rect 47075 31297 47084 31331
rect 47032 31288 47084 31297
rect 4712 31084 4764 31136
rect 46940 31127 46992 31136
rect 46940 31093 46949 31127
rect 46949 31093 46983 31127
rect 46983 31093 46992 31127
rect 46940 31084 46992 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 48412 30787 48464 30796
rect 48412 30753 48421 30787
rect 48421 30753 48455 30787
rect 48455 30753 48464 30787
rect 49240 30787 49292 30796
rect 48412 30744 48464 30753
rect 49240 30753 49249 30787
rect 49249 30753 49283 30787
rect 49283 30753 49292 30787
rect 49240 30744 49292 30753
rect 46296 30719 46348 30728
rect 46296 30685 46305 30719
rect 46305 30685 46339 30719
rect 46339 30685 46348 30719
rect 46296 30676 46348 30685
rect 46940 30719 46992 30728
rect 46940 30685 46949 30719
rect 46949 30685 46983 30719
rect 46983 30685 46992 30719
rect 46940 30676 46992 30685
rect 48320 30676 48372 30728
rect 58164 30676 58216 30728
rect 2412 30608 2464 30660
rect 58256 30583 58308 30592
rect 58256 30549 58265 30583
rect 58265 30549 58299 30583
rect 58299 30549 58308 30583
rect 58256 30540 58308 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 46756 30336 46808 30388
rect 44824 30311 44876 30320
rect 44824 30277 44833 30311
rect 44833 30277 44867 30311
rect 44867 30277 44876 30311
rect 44824 30268 44876 30277
rect 46296 30268 46348 30320
rect 48320 30268 48372 30320
rect 49516 30268 49568 30320
rect 46388 30243 46440 30252
rect 46388 30209 46397 30243
rect 46397 30209 46431 30243
rect 46431 30209 46440 30243
rect 46388 30200 46440 30209
rect 49240 30200 49292 30252
rect 44916 30064 44968 30116
rect 49424 30039 49476 30048
rect 49424 30005 49433 30039
rect 49433 30005 49467 30039
rect 49467 30005 49476 30039
rect 49424 29996 49476 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 46756 29835 46808 29844
rect 46756 29801 46765 29835
rect 46765 29801 46799 29835
rect 46799 29801 46808 29835
rect 46756 29792 46808 29801
rect 47032 29792 47084 29844
rect 48412 29792 48464 29844
rect 46388 29724 46440 29776
rect 48136 29767 48188 29776
rect 44732 29656 44784 29708
rect 46112 29656 46164 29708
rect 45468 29588 45520 29640
rect 46204 29588 46256 29640
rect 48136 29733 48145 29767
rect 48145 29733 48179 29767
rect 48179 29733 48188 29767
rect 48136 29724 48188 29733
rect 48964 29767 49016 29776
rect 48964 29733 48973 29767
rect 48973 29733 49007 29767
rect 49007 29733 49016 29767
rect 48964 29724 49016 29733
rect 57520 29724 57572 29776
rect 49240 29699 49292 29708
rect 49240 29665 49249 29699
rect 49249 29665 49283 29699
rect 49283 29665 49292 29699
rect 49240 29656 49292 29665
rect 50988 29631 51040 29640
rect 47952 29520 48004 29572
rect 50988 29597 50997 29631
rect 50997 29597 51031 29631
rect 51031 29597 51040 29631
rect 50988 29588 51040 29597
rect 51816 29588 51868 29640
rect 1676 29495 1728 29504
rect 1676 29461 1685 29495
rect 1685 29461 1719 29495
rect 1719 29461 1728 29495
rect 1676 29452 1728 29461
rect 2412 29495 2464 29504
rect 2412 29461 2421 29495
rect 2421 29461 2455 29495
rect 2455 29461 2464 29495
rect 2412 29452 2464 29461
rect 45192 29495 45244 29504
rect 45192 29461 45201 29495
rect 45201 29461 45235 29495
rect 45235 29461 45244 29495
rect 45192 29452 45244 29461
rect 47216 29452 47268 29504
rect 50988 29452 51040 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 44824 29248 44876 29300
rect 46112 29291 46164 29300
rect 46112 29257 46137 29291
rect 46137 29257 46164 29291
rect 46112 29248 46164 29257
rect 46388 29248 46440 29300
rect 49608 29248 49660 29300
rect 51816 29291 51868 29300
rect 44824 29112 44876 29164
rect 45468 29112 45520 29164
rect 47216 29112 47268 29164
rect 47952 29155 48004 29164
rect 47952 29121 47961 29155
rect 47961 29121 47995 29155
rect 47995 29121 48004 29155
rect 47952 29112 48004 29121
rect 49240 29155 49292 29164
rect 49240 29121 49249 29155
rect 49249 29121 49283 29155
rect 49283 29121 49292 29155
rect 49240 29112 49292 29121
rect 49516 29112 49568 29164
rect 49792 29112 49844 29164
rect 51816 29257 51825 29291
rect 51825 29257 51859 29291
rect 51859 29257 51868 29291
rect 51816 29248 51868 29257
rect 50896 29180 50948 29232
rect 44732 29087 44784 29096
rect 44732 29053 44741 29087
rect 44741 29053 44775 29087
rect 44775 29053 44784 29087
rect 44732 29044 44784 29053
rect 48964 29044 49016 29096
rect 49332 29044 49384 29096
rect 51172 29112 51224 29164
rect 54116 29112 54168 29164
rect 55220 29112 55272 29164
rect 1860 28976 1912 29028
rect 46204 28908 46256 28960
rect 46848 28951 46900 28960
rect 46848 28917 46857 28951
rect 46857 28917 46891 28951
rect 46891 28917 46900 28951
rect 46848 28908 46900 28917
rect 48136 28951 48188 28960
rect 48136 28917 48145 28951
rect 48145 28917 48179 28951
rect 48179 28917 48188 28951
rect 48136 28908 48188 28917
rect 50988 28951 51040 28960
rect 50988 28917 50997 28951
rect 50997 28917 51031 28951
rect 51031 28917 51040 28951
rect 50988 28908 51040 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 46204 28747 46256 28756
rect 46204 28713 46213 28747
rect 46213 28713 46247 28747
rect 46247 28713 46256 28747
rect 46204 28704 46256 28713
rect 47216 28747 47268 28756
rect 46020 28636 46072 28688
rect 47216 28713 47225 28747
rect 47225 28713 47259 28747
rect 47259 28713 47268 28747
rect 47216 28704 47268 28713
rect 46848 28611 46900 28620
rect 46848 28577 46857 28611
rect 46857 28577 46891 28611
rect 46891 28577 46900 28611
rect 46848 28568 46900 28577
rect 45652 28500 45704 28552
rect 49332 28568 49384 28620
rect 45008 28432 45060 28484
rect 49424 28543 49476 28552
rect 45652 28364 45704 28416
rect 46664 28364 46716 28416
rect 49424 28509 49433 28543
rect 49433 28509 49467 28543
rect 49467 28509 49476 28543
rect 49424 28500 49476 28509
rect 49608 28543 49660 28552
rect 49608 28509 49617 28543
rect 49617 28509 49651 28543
rect 49651 28509 49660 28543
rect 49608 28500 49660 28509
rect 50804 28636 50856 28688
rect 50988 28568 51040 28620
rect 51356 28543 51408 28552
rect 51356 28509 51365 28543
rect 51365 28509 51399 28543
rect 51399 28509 51408 28543
rect 51356 28500 51408 28509
rect 52920 28543 52972 28552
rect 49792 28432 49844 28484
rect 51172 28432 51224 28484
rect 52920 28509 52929 28543
rect 52929 28509 52963 28543
rect 52963 28509 52972 28543
rect 52920 28500 52972 28509
rect 53932 28568 53984 28620
rect 53748 28500 53800 28552
rect 57152 28500 57204 28552
rect 57244 28432 57296 28484
rect 50068 28364 50120 28416
rect 53012 28407 53064 28416
rect 53012 28373 53021 28407
rect 53021 28373 53055 28407
rect 53055 28373 53064 28407
rect 53012 28364 53064 28373
rect 53840 28407 53892 28416
rect 53840 28373 53849 28407
rect 53849 28373 53883 28407
rect 53883 28373 53892 28407
rect 53840 28364 53892 28373
rect 56968 28407 57020 28416
rect 56968 28373 56977 28407
rect 56977 28373 57011 28407
rect 57011 28373 57020 28407
rect 56968 28364 57020 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 46848 28160 46900 28212
rect 2504 28092 2556 28144
rect 45744 28092 45796 28144
rect 57244 28092 57296 28144
rect 44640 28067 44692 28076
rect 44640 28033 44649 28067
rect 44649 28033 44683 28067
rect 44683 28033 44692 28067
rect 44640 28024 44692 28033
rect 45100 28067 45152 28076
rect 45100 28033 45109 28067
rect 45109 28033 45143 28067
rect 45143 28033 45152 28067
rect 45100 28024 45152 28033
rect 45836 28024 45888 28076
rect 47860 28067 47912 28076
rect 46296 27956 46348 28008
rect 47860 28033 47869 28067
rect 47869 28033 47903 28067
rect 47903 28033 47912 28067
rect 47860 28024 47912 28033
rect 48504 28067 48556 28076
rect 47492 27956 47544 28008
rect 48504 28033 48513 28067
rect 48513 28033 48547 28067
rect 48547 28033 48556 28067
rect 48504 28024 48556 28033
rect 49700 28067 49752 28076
rect 49700 28033 49709 28067
rect 49709 28033 49743 28067
rect 49743 28033 49752 28067
rect 49700 28024 49752 28033
rect 50620 28024 50672 28076
rect 49424 27956 49476 28008
rect 49792 27999 49844 28008
rect 49792 27965 49801 27999
rect 49801 27965 49835 27999
rect 49835 27965 49844 27999
rect 50804 28024 50856 28076
rect 51356 28067 51408 28076
rect 51356 28033 51365 28067
rect 51365 28033 51399 28067
rect 51399 28033 51408 28067
rect 51356 28024 51408 28033
rect 51080 27999 51132 28008
rect 49792 27956 49844 27965
rect 51080 27965 51089 27999
rect 51089 27965 51123 27999
rect 51123 27965 51132 27999
rect 51080 27956 51132 27965
rect 52828 28024 52880 28076
rect 53012 28024 53064 28076
rect 53748 28024 53800 28076
rect 54208 28024 54260 28076
rect 54392 28067 54444 28076
rect 54392 28033 54401 28067
rect 54401 28033 54435 28067
rect 54435 28033 54444 28067
rect 54392 28024 54444 28033
rect 55588 28024 55640 28076
rect 55864 28067 55916 28076
rect 55864 28033 55873 28067
rect 55873 28033 55907 28067
rect 55907 28033 55916 28067
rect 55864 28024 55916 28033
rect 56048 28024 56100 28076
rect 45928 27888 45980 27940
rect 50988 27888 51040 27940
rect 53932 27956 53984 28008
rect 55220 27999 55272 28008
rect 55220 27965 55229 27999
rect 55229 27965 55263 27999
rect 55263 27965 55272 27999
rect 55220 27956 55272 27965
rect 47124 27863 47176 27872
rect 47124 27829 47133 27863
rect 47133 27829 47167 27863
rect 47167 27829 47176 27863
rect 47124 27820 47176 27829
rect 53196 27820 53248 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 46020 27616 46072 27668
rect 47216 27659 47268 27668
rect 47216 27625 47225 27659
rect 47225 27625 47259 27659
rect 47259 27625 47268 27659
rect 47216 27616 47268 27625
rect 49608 27616 49660 27668
rect 51356 27616 51408 27668
rect 45652 27548 45704 27600
rect 47860 27548 47912 27600
rect 47952 27548 48004 27600
rect 54208 27548 54260 27600
rect 55588 27591 55640 27600
rect 55588 27557 55597 27591
rect 55597 27557 55631 27591
rect 55631 27557 55640 27591
rect 55588 27548 55640 27557
rect 44640 27523 44692 27532
rect 44640 27489 44649 27523
rect 44649 27489 44683 27523
rect 44683 27489 44692 27523
rect 44640 27480 44692 27489
rect 45928 27523 45980 27532
rect 43904 27455 43956 27464
rect 43904 27421 43913 27455
rect 43913 27421 43947 27455
rect 43947 27421 43956 27455
rect 43904 27412 43956 27421
rect 43996 27455 44048 27464
rect 43996 27421 44005 27455
rect 44005 27421 44039 27455
rect 44039 27421 44048 27455
rect 44180 27455 44232 27464
rect 43996 27412 44048 27421
rect 44180 27421 44189 27455
rect 44189 27421 44223 27455
rect 44223 27421 44232 27455
rect 44180 27412 44232 27421
rect 44456 27412 44508 27464
rect 45928 27489 45937 27523
rect 45937 27489 45971 27523
rect 45971 27489 45980 27523
rect 45928 27480 45980 27489
rect 47492 27480 47544 27532
rect 45744 27455 45796 27464
rect 45744 27421 45753 27455
rect 45753 27421 45787 27455
rect 45787 27421 45796 27455
rect 45744 27412 45796 27421
rect 45836 27455 45888 27464
rect 45836 27421 45845 27455
rect 45845 27421 45879 27455
rect 45879 27421 45888 27455
rect 45836 27412 45888 27421
rect 46296 27412 46348 27464
rect 46664 27412 46716 27464
rect 47308 27412 47360 27464
rect 52276 27523 52328 27532
rect 52276 27489 52285 27523
rect 52285 27489 52319 27523
rect 52319 27489 52328 27523
rect 52276 27480 52328 27489
rect 52920 27523 52972 27532
rect 52920 27489 52929 27523
rect 52929 27489 52963 27523
rect 52963 27489 52972 27523
rect 52920 27480 52972 27489
rect 49424 27455 49476 27464
rect 49424 27421 49433 27455
rect 49433 27421 49467 27455
rect 49467 27421 49476 27455
rect 49424 27412 49476 27421
rect 49700 27455 49752 27464
rect 49700 27421 49709 27455
rect 49709 27421 49743 27455
rect 49743 27421 49752 27455
rect 49700 27412 49752 27421
rect 50620 27455 50672 27464
rect 50620 27421 50629 27455
rect 50629 27421 50663 27455
rect 50663 27421 50672 27455
rect 50620 27412 50672 27421
rect 50896 27455 50948 27464
rect 50896 27421 50905 27455
rect 50905 27421 50939 27455
rect 50939 27421 50948 27455
rect 50896 27412 50948 27421
rect 52368 27455 52420 27464
rect 52368 27421 52377 27455
rect 52377 27421 52411 27455
rect 52411 27421 52420 27455
rect 52368 27412 52420 27421
rect 54392 27480 54444 27532
rect 53748 27412 53800 27464
rect 53932 27455 53984 27464
rect 53932 27421 53941 27455
rect 53941 27421 53975 27455
rect 53975 27421 53984 27455
rect 54116 27455 54168 27464
rect 53932 27412 53984 27421
rect 54116 27421 54125 27455
rect 54125 27421 54159 27455
rect 54159 27421 54168 27455
rect 54116 27412 54168 27421
rect 54576 27455 54628 27464
rect 54576 27421 54585 27455
rect 54585 27421 54619 27455
rect 54619 27421 54628 27455
rect 54576 27412 54628 27421
rect 55220 27412 55272 27464
rect 56968 27455 57020 27464
rect 56968 27421 56977 27455
rect 56977 27421 57011 27455
rect 57011 27421 57020 27455
rect 56968 27412 57020 27421
rect 57888 27455 57940 27464
rect 57888 27421 57897 27455
rect 57897 27421 57931 27455
rect 57931 27421 57940 27455
rect 57888 27412 57940 27421
rect 2412 27344 2464 27396
rect 49516 27276 49568 27328
rect 50712 27319 50764 27328
rect 50712 27285 50721 27319
rect 50721 27285 50755 27319
rect 50755 27285 50764 27319
rect 50712 27276 50764 27285
rect 53932 27276 53984 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 45744 27072 45796 27124
rect 47308 27072 47360 27124
rect 48504 27072 48556 27124
rect 51172 27115 51224 27124
rect 51172 27081 51181 27115
rect 51181 27081 51215 27115
rect 51215 27081 51224 27115
rect 51172 27072 51224 27081
rect 54392 27115 54444 27124
rect 44456 27004 44508 27056
rect 43812 26936 43864 26988
rect 43904 26936 43956 26988
rect 44640 26936 44692 26988
rect 12440 26800 12492 26852
rect 44272 26868 44324 26920
rect 44916 26911 44968 26920
rect 44916 26877 44925 26911
rect 44925 26877 44959 26911
rect 44959 26877 44968 26911
rect 44916 26868 44968 26877
rect 47124 27004 47176 27056
rect 47584 27004 47636 27056
rect 50712 27004 50764 27056
rect 50896 27004 50948 27056
rect 53012 27004 53064 27056
rect 54392 27081 54401 27115
rect 54401 27081 54435 27115
rect 54435 27081 54444 27115
rect 54392 27072 54444 27081
rect 57152 27072 57204 27124
rect 54576 27004 54628 27056
rect 46572 26936 46624 26988
rect 48044 26979 48096 26988
rect 48044 26945 48053 26979
rect 48053 26945 48087 26979
rect 48087 26945 48096 26979
rect 48044 26936 48096 26945
rect 48136 26979 48188 26988
rect 48136 26945 48145 26979
rect 48145 26945 48179 26979
rect 48179 26945 48188 26979
rect 48136 26936 48188 26945
rect 49240 26936 49292 26988
rect 52276 26936 52328 26988
rect 52368 26979 52420 26988
rect 52368 26945 52377 26979
rect 52377 26945 52411 26979
rect 52411 26945 52420 26979
rect 54300 26979 54352 26988
rect 52368 26936 52420 26945
rect 54300 26945 54309 26979
rect 54309 26945 54343 26979
rect 54343 26945 54352 26979
rect 54300 26936 54352 26945
rect 54944 26936 54996 26988
rect 55864 26979 55916 26988
rect 46020 26868 46072 26920
rect 47952 26868 48004 26920
rect 55864 26945 55873 26979
rect 55873 26945 55907 26979
rect 55907 26945 55916 26979
rect 55864 26936 55916 26945
rect 56048 26979 56100 26988
rect 56048 26945 56057 26979
rect 56057 26945 56091 26979
rect 56091 26945 56100 26979
rect 56048 26936 56100 26945
rect 56968 26936 57020 26988
rect 56324 26868 56376 26920
rect 57244 26911 57296 26920
rect 57244 26877 57253 26911
rect 57253 26877 57287 26911
rect 57287 26877 57296 26911
rect 57244 26868 57296 26877
rect 44180 26800 44232 26852
rect 48228 26800 48280 26852
rect 53196 26843 53248 26852
rect 53196 26809 53205 26843
rect 53205 26809 53239 26843
rect 53239 26809 53248 26843
rect 53196 26800 53248 26809
rect 57060 26800 57112 26852
rect 44916 26732 44968 26784
rect 45100 26732 45152 26784
rect 46112 26775 46164 26784
rect 46112 26741 46121 26775
rect 46121 26741 46155 26775
rect 46155 26741 46164 26775
rect 46112 26732 46164 26741
rect 46664 26732 46716 26784
rect 48780 26732 48832 26784
rect 50620 26732 50672 26784
rect 53380 26775 53432 26784
rect 53380 26741 53389 26775
rect 53389 26741 53423 26775
rect 53423 26741 53432 26775
rect 53380 26732 53432 26741
rect 55220 26775 55272 26784
rect 55220 26741 55229 26775
rect 55229 26741 55263 26775
rect 55263 26741 55272 26775
rect 57520 26775 57572 26784
rect 55220 26732 55272 26741
rect 57520 26741 57529 26775
rect 57529 26741 57563 26775
rect 57563 26741 57572 26775
rect 57520 26732 57572 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 43904 26528 43956 26580
rect 40040 26460 40092 26512
rect 43812 26460 43864 26512
rect 46112 26528 46164 26580
rect 47032 26571 47084 26580
rect 47032 26537 47041 26571
rect 47041 26537 47075 26571
rect 47075 26537 47084 26571
rect 47032 26528 47084 26537
rect 47216 26528 47268 26580
rect 49700 26528 49752 26580
rect 50988 26528 51040 26580
rect 53380 26528 53432 26580
rect 58532 26528 58584 26580
rect 45928 26460 45980 26512
rect 46204 26460 46256 26512
rect 46572 26392 46624 26444
rect 48044 26460 48096 26512
rect 47952 26435 48004 26444
rect 47952 26401 47961 26435
rect 47961 26401 47995 26435
rect 47995 26401 48004 26435
rect 47952 26392 48004 26401
rect 45376 26367 45428 26376
rect 45376 26333 45385 26367
rect 45385 26333 45419 26367
rect 45419 26333 45428 26367
rect 45376 26324 45428 26333
rect 46020 26324 46072 26376
rect 46940 26367 46992 26376
rect 38476 26299 38528 26308
rect 38476 26265 38485 26299
rect 38485 26265 38519 26299
rect 38519 26265 38528 26299
rect 38476 26256 38528 26265
rect 44272 26299 44324 26308
rect 44272 26265 44299 26299
rect 44299 26265 44324 26299
rect 44272 26256 44324 26265
rect 44456 26299 44508 26308
rect 44456 26265 44465 26299
rect 44465 26265 44499 26299
rect 44499 26265 44508 26299
rect 44456 26256 44508 26265
rect 45836 26256 45888 26308
rect 46940 26333 46949 26367
rect 46949 26333 46983 26367
rect 46983 26333 46992 26367
rect 46940 26324 46992 26333
rect 47584 26324 47636 26376
rect 48228 26460 48280 26512
rect 54944 26460 54996 26512
rect 56508 26460 56560 26512
rect 56968 26460 57020 26512
rect 57428 26460 57480 26512
rect 57888 26435 57940 26444
rect 57888 26401 57897 26435
rect 57897 26401 57931 26435
rect 57931 26401 57940 26435
rect 57888 26392 57940 26401
rect 48780 26367 48832 26376
rect 48780 26333 48789 26367
rect 48789 26333 48823 26367
rect 48823 26333 48832 26367
rect 48780 26324 48832 26333
rect 49148 26367 49200 26376
rect 49148 26333 49157 26367
rect 49157 26333 49191 26367
rect 49191 26333 49200 26367
rect 49148 26324 49200 26333
rect 49240 26367 49292 26376
rect 49240 26333 49249 26367
rect 49249 26333 49283 26367
rect 49283 26333 49292 26367
rect 49240 26324 49292 26333
rect 49516 26324 49568 26376
rect 50620 26367 50672 26376
rect 50620 26333 50629 26367
rect 50629 26333 50663 26367
rect 50663 26333 50672 26367
rect 50620 26324 50672 26333
rect 50712 26367 50764 26376
rect 50712 26333 50721 26367
rect 50721 26333 50755 26367
rect 50755 26333 50764 26367
rect 53840 26367 53892 26376
rect 50712 26324 50764 26333
rect 53840 26333 53849 26367
rect 53849 26333 53883 26367
rect 53883 26333 53892 26367
rect 53840 26324 53892 26333
rect 54024 26367 54076 26376
rect 54024 26333 54033 26367
rect 54033 26333 54067 26367
rect 54067 26333 54076 26367
rect 54024 26324 54076 26333
rect 56324 26324 56376 26376
rect 56508 26367 56560 26376
rect 56508 26333 56517 26367
rect 56517 26333 56551 26367
rect 56551 26333 56560 26367
rect 56508 26324 56560 26333
rect 58256 26367 58308 26376
rect 58256 26333 58265 26367
rect 58265 26333 58299 26367
rect 58299 26333 58308 26367
rect 58256 26324 58308 26333
rect 38936 26231 38988 26240
rect 38936 26197 38945 26231
rect 38945 26197 38979 26231
rect 38979 26197 38988 26231
rect 38936 26188 38988 26197
rect 47124 26256 47176 26308
rect 48044 26299 48096 26308
rect 48044 26265 48053 26299
rect 48053 26265 48087 26299
rect 48087 26265 48096 26299
rect 48044 26256 48096 26265
rect 49608 26299 49660 26308
rect 49608 26265 49617 26299
rect 49617 26265 49651 26299
rect 49651 26265 49660 26299
rect 49608 26256 49660 26265
rect 50804 26256 50856 26308
rect 55956 26256 56008 26308
rect 57060 26256 57112 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 44732 25984 44784 26036
rect 44272 25916 44324 25968
rect 38936 25891 38988 25900
rect 38936 25857 38945 25891
rect 38945 25857 38979 25891
rect 38979 25857 38988 25891
rect 38936 25848 38988 25857
rect 39028 25891 39080 25900
rect 39028 25857 39037 25891
rect 39037 25857 39071 25891
rect 39071 25857 39080 25891
rect 39028 25848 39080 25857
rect 44732 25848 44784 25900
rect 45376 25916 45428 25968
rect 45744 25959 45796 25968
rect 45744 25925 45753 25959
rect 45753 25925 45787 25959
rect 45787 25925 45796 25959
rect 45744 25916 45796 25925
rect 43904 25823 43956 25832
rect 43904 25789 43913 25823
rect 43913 25789 43947 25823
rect 43947 25789 43956 25823
rect 43904 25780 43956 25789
rect 46572 25891 46624 25900
rect 46572 25857 46581 25891
rect 46581 25857 46615 25891
rect 46615 25857 46624 25891
rect 46572 25848 46624 25857
rect 48044 25984 48096 26036
rect 54024 26027 54076 26036
rect 54024 25993 54033 26027
rect 54033 25993 54067 26027
rect 54067 25993 54076 26027
rect 54024 25984 54076 25993
rect 57152 25984 57204 26036
rect 48780 25916 48832 25968
rect 49608 25916 49660 25968
rect 46940 25848 46992 25900
rect 48872 25848 48924 25900
rect 49424 25891 49476 25900
rect 49424 25857 49433 25891
rect 49433 25857 49467 25891
rect 49467 25857 49476 25891
rect 49424 25848 49476 25857
rect 49884 25848 49936 25900
rect 50712 25891 50764 25900
rect 50712 25857 50721 25891
rect 50721 25857 50755 25891
rect 50755 25857 50764 25891
rect 50712 25848 50764 25857
rect 50988 25891 51040 25900
rect 50988 25857 50997 25891
rect 50997 25857 51031 25891
rect 51031 25857 51040 25891
rect 50988 25848 51040 25857
rect 53196 25848 53248 25900
rect 46112 25780 46164 25832
rect 47032 25780 47084 25832
rect 49240 25823 49292 25832
rect 49240 25789 49249 25823
rect 49249 25789 49283 25823
rect 49283 25789 49292 25823
rect 49240 25780 49292 25789
rect 52184 25780 52236 25832
rect 52736 25780 52788 25832
rect 54300 25848 54352 25900
rect 54392 25848 54444 25900
rect 55036 25891 55088 25900
rect 55036 25857 55045 25891
rect 55045 25857 55079 25891
rect 55079 25857 55088 25891
rect 56048 25891 56100 25900
rect 55036 25848 55088 25857
rect 56048 25857 56057 25891
rect 56057 25857 56091 25891
rect 56091 25857 56100 25891
rect 56048 25848 56100 25857
rect 57060 25891 57112 25900
rect 57060 25857 57069 25891
rect 57069 25857 57103 25891
rect 57103 25857 57112 25891
rect 57060 25848 57112 25857
rect 57152 25891 57204 25900
rect 57152 25857 57161 25891
rect 57161 25857 57195 25891
rect 57195 25857 57204 25891
rect 57428 25891 57480 25900
rect 57152 25848 57204 25857
rect 57428 25857 57437 25891
rect 57437 25857 57471 25891
rect 57471 25857 57480 25891
rect 57428 25848 57480 25857
rect 57612 25848 57664 25900
rect 55864 25780 55916 25832
rect 58256 25848 58308 25900
rect 47124 25712 47176 25764
rect 49516 25712 49568 25764
rect 54208 25712 54260 25764
rect 1952 25644 2004 25696
rect 46020 25644 46072 25696
rect 47676 25644 47728 25696
rect 49148 25687 49200 25696
rect 49148 25653 49157 25687
rect 49157 25653 49191 25687
rect 49191 25653 49200 25687
rect 49148 25644 49200 25653
rect 52460 25644 52512 25696
rect 53288 25687 53340 25696
rect 53288 25653 53297 25687
rect 53297 25653 53331 25687
rect 53331 25653 53340 25687
rect 53288 25644 53340 25653
rect 55220 25644 55272 25696
rect 55956 25644 56008 25696
rect 56876 25687 56928 25696
rect 56876 25653 56885 25687
rect 56885 25653 56919 25687
rect 56919 25653 56928 25687
rect 56876 25644 56928 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 40408 25483 40460 25492
rect 40408 25449 40417 25483
rect 40417 25449 40451 25483
rect 40451 25449 40460 25483
rect 40408 25440 40460 25449
rect 43904 25483 43956 25492
rect 43904 25449 43913 25483
rect 43913 25449 43947 25483
rect 43947 25449 43956 25483
rect 43904 25440 43956 25449
rect 45192 25440 45244 25492
rect 46020 25440 46072 25492
rect 47492 25483 47544 25492
rect 47492 25449 47501 25483
rect 47501 25449 47535 25483
rect 47535 25449 47544 25483
rect 47492 25440 47544 25449
rect 48780 25483 48832 25492
rect 48780 25449 48789 25483
rect 48789 25449 48823 25483
rect 48823 25449 48832 25483
rect 48780 25440 48832 25449
rect 50804 25483 50856 25492
rect 50804 25449 50813 25483
rect 50813 25449 50847 25483
rect 50847 25449 50856 25483
rect 50804 25440 50856 25449
rect 54300 25440 54352 25492
rect 55956 25483 56008 25492
rect 55956 25449 55965 25483
rect 55965 25449 55999 25483
rect 55999 25449 56008 25483
rect 55956 25440 56008 25449
rect 57060 25440 57112 25492
rect 57796 25440 57848 25492
rect 57612 25372 57664 25424
rect 39028 25304 39080 25356
rect 44456 25304 44508 25356
rect 46204 25304 46256 25356
rect 47308 25347 47360 25356
rect 47308 25313 47317 25347
rect 47317 25313 47351 25347
rect 47351 25313 47360 25347
rect 47308 25304 47360 25313
rect 50712 25304 50764 25356
rect 52368 25304 52420 25356
rect 52828 25347 52880 25356
rect 52828 25313 52837 25347
rect 52837 25313 52871 25347
rect 52871 25313 52880 25347
rect 52828 25304 52880 25313
rect 54392 25304 54444 25356
rect 56140 25347 56192 25356
rect 56140 25313 56149 25347
rect 56149 25313 56183 25347
rect 56183 25313 56192 25347
rect 56140 25304 56192 25313
rect 37740 25236 37792 25288
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 38200 25279 38252 25288
rect 38200 25245 38209 25279
rect 38209 25245 38243 25279
rect 38243 25245 38252 25279
rect 38200 25236 38252 25245
rect 38844 25279 38896 25288
rect 38844 25245 38853 25279
rect 38853 25245 38887 25279
rect 38887 25245 38896 25279
rect 38844 25236 38896 25245
rect 39212 25279 39264 25288
rect 39212 25245 39221 25279
rect 39221 25245 39255 25279
rect 39255 25245 39264 25279
rect 39212 25236 39264 25245
rect 39396 25279 39448 25288
rect 39396 25245 39405 25279
rect 39405 25245 39439 25279
rect 39439 25245 39448 25279
rect 39396 25236 39448 25245
rect 40040 25279 40092 25288
rect 40040 25245 40049 25279
rect 40049 25245 40083 25279
rect 40083 25245 40092 25279
rect 40040 25236 40092 25245
rect 40224 25279 40276 25288
rect 40224 25245 40233 25279
rect 40233 25245 40267 25279
rect 40267 25245 40276 25279
rect 40224 25236 40276 25245
rect 37188 25211 37240 25220
rect 37188 25177 37197 25211
rect 37197 25177 37231 25211
rect 37231 25177 37240 25211
rect 37188 25168 37240 25177
rect 44916 25236 44968 25288
rect 45836 25236 45888 25288
rect 48504 25279 48556 25288
rect 37464 25100 37516 25152
rect 44088 25100 44140 25152
rect 47124 25168 47176 25220
rect 45468 25100 45520 25152
rect 45652 25143 45704 25152
rect 45652 25109 45661 25143
rect 45661 25109 45695 25143
rect 45695 25109 45704 25143
rect 48504 25245 48513 25279
rect 48513 25245 48547 25279
rect 48547 25245 48556 25279
rect 48504 25236 48556 25245
rect 49516 25279 49568 25288
rect 49516 25245 49525 25279
rect 49525 25245 49559 25279
rect 49559 25245 49568 25279
rect 49516 25236 49568 25245
rect 48964 25168 49016 25220
rect 50988 25236 51040 25288
rect 53288 25236 53340 25288
rect 53932 25279 53984 25288
rect 53932 25245 53941 25279
rect 53941 25245 53975 25279
rect 53975 25245 53984 25279
rect 53932 25236 53984 25245
rect 54208 25236 54260 25288
rect 55036 25236 55088 25288
rect 55864 25279 55916 25288
rect 55864 25245 55873 25279
rect 55873 25245 55907 25279
rect 55907 25245 55916 25279
rect 55864 25236 55916 25245
rect 57520 25236 57572 25288
rect 57060 25168 57112 25220
rect 45652 25100 45704 25109
rect 49792 25100 49844 25152
rect 58440 25100 58492 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 37188 24896 37240 24948
rect 38200 24896 38252 24948
rect 40224 24939 40276 24948
rect 37464 24871 37516 24880
rect 37464 24837 37473 24871
rect 37473 24837 37507 24871
rect 37507 24837 37516 24871
rect 37464 24828 37516 24837
rect 35348 24760 35400 24812
rect 36452 24760 36504 24812
rect 38384 24760 38436 24812
rect 40224 24905 40233 24939
rect 40233 24905 40267 24939
rect 40267 24905 40276 24939
rect 40224 24896 40276 24905
rect 47308 24896 47360 24948
rect 48504 24896 48556 24948
rect 49424 24896 49476 24948
rect 44916 24828 44968 24880
rect 31668 24692 31720 24744
rect 34796 24692 34848 24744
rect 36360 24692 36412 24744
rect 39948 24760 40000 24812
rect 40316 24803 40368 24812
rect 40316 24769 40325 24803
rect 40325 24769 40359 24803
rect 40359 24769 40368 24803
rect 40316 24760 40368 24769
rect 43812 24803 43864 24812
rect 43812 24769 43821 24803
rect 43821 24769 43855 24803
rect 43855 24769 43864 24803
rect 43812 24760 43864 24769
rect 45468 24760 45520 24812
rect 47124 24828 47176 24880
rect 46204 24760 46256 24812
rect 46572 24760 46624 24812
rect 49792 24828 49844 24880
rect 50988 24896 51040 24948
rect 40040 24692 40092 24744
rect 45560 24735 45612 24744
rect 45560 24701 45569 24735
rect 45569 24701 45603 24735
rect 45603 24701 45612 24735
rect 45560 24692 45612 24701
rect 45836 24735 45888 24744
rect 45836 24701 45845 24735
rect 45845 24701 45879 24735
rect 45879 24701 45888 24735
rect 45836 24692 45888 24701
rect 46020 24692 46072 24744
rect 35624 24624 35676 24676
rect 38844 24624 38896 24676
rect 39396 24624 39448 24676
rect 44272 24667 44324 24676
rect 44272 24633 44281 24667
rect 44281 24633 44315 24667
rect 44315 24633 44324 24667
rect 44272 24624 44324 24633
rect 49516 24760 49568 24812
rect 49884 24760 49936 24812
rect 52736 24828 52788 24880
rect 52460 24760 52512 24812
rect 52920 24803 52972 24812
rect 52920 24769 52929 24803
rect 52929 24769 52963 24803
rect 52963 24769 52972 24803
rect 52920 24760 52972 24769
rect 53196 24803 53248 24812
rect 49976 24692 50028 24744
rect 53196 24769 53205 24803
rect 53205 24769 53239 24803
rect 53239 24769 53248 24803
rect 53196 24760 53248 24769
rect 53932 24760 53984 24812
rect 54760 24803 54812 24812
rect 54760 24769 54769 24803
rect 54769 24769 54803 24803
rect 54803 24769 54812 24803
rect 54760 24760 54812 24769
rect 55496 24803 55548 24812
rect 55496 24769 55505 24803
rect 55505 24769 55539 24803
rect 55539 24769 55548 24803
rect 55496 24760 55548 24769
rect 56324 24760 56376 24812
rect 56416 24735 56468 24744
rect 56416 24701 56425 24735
rect 56425 24701 56459 24735
rect 56459 24701 56468 24735
rect 56416 24692 56468 24701
rect 56508 24692 56560 24744
rect 58440 24760 58492 24812
rect 37740 24556 37792 24608
rect 43904 24556 43956 24608
rect 44732 24556 44784 24608
rect 45376 24599 45428 24608
rect 45376 24565 45385 24599
rect 45385 24565 45419 24599
rect 45419 24565 45428 24599
rect 45376 24556 45428 24565
rect 45744 24556 45796 24608
rect 50068 24624 50120 24676
rect 48964 24599 49016 24608
rect 48964 24565 48973 24599
rect 48973 24565 49007 24599
rect 49007 24565 49016 24599
rect 48964 24556 49016 24565
rect 50160 24599 50212 24608
rect 50160 24565 50169 24599
rect 50169 24565 50203 24599
rect 50203 24565 50212 24599
rect 50160 24556 50212 24565
rect 56968 24556 57020 24608
rect 58256 24599 58308 24608
rect 58256 24565 58265 24599
rect 58265 24565 58299 24599
rect 58299 24565 58308 24599
rect 58256 24556 58308 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 35624 24352 35676 24404
rect 36268 24352 36320 24404
rect 37464 24352 37516 24404
rect 38384 24395 38436 24404
rect 38384 24361 38393 24395
rect 38393 24361 38427 24395
rect 38427 24361 38436 24395
rect 38384 24352 38436 24361
rect 40040 24395 40092 24404
rect 40040 24361 40049 24395
rect 40049 24361 40083 24395
rect 40083 24361 40092 24395
rect 40040 24352 40092 24361
rect 43996 24395 44048 24404
rect 43996 24361 44005 24395
rect 44005 24361 44039 24395
rect 44039 24361 44048 24395
rect 43996 24352 44048 24361
rect 45192 24352 45244 24404
rect 47124 24352 47176 24404
rect 50712 24352 50764 24404
rect 55864 24395 55916 24404
rect 55864 24361 55873 24395
rect 55873 24361 55907 24395
rect 55907 24361 55916 24395
rect 55864 24352 55916 24361
rect 58072 24352 58124 24404
rect 43904 24284 43956 24336
rect 34796 24216 34848 24268
rect 38752 24216 38804 24268
rect 40316 24216 40368 24268
rect 27068 24148 27120 24200
rect 27620 24148 27672 24200
rect 31484 24148 31536 24200
rect 31576 24148 31628 24200
rect 32496 24191 32548 24200
rect 32496 24157 32505 24191
rect 32505 24157 32539 24191
rect 32539 24157 32548 24191
rect 32496 24148 32548 24157
rect 35256 24191 35308 24200
rect 35256 24157 35265 24191
rect 35265 24157 35299 24191
rect 35299 24157 35308 24191
rect 35256 24148 35308 24157
rect 36452 24148 36504 24200
rect 38016 24148 38068 24200
rect 38476 24148 38528 24200
rect 40132 24148 40184 24200
rect 40592 24191 40644 24200
rect 40592 24157 40601 24191
rect 40601 24157 40635 24191
rect 40635 24157 40644 24191
rect 40592 24148 40644 24157
rect 10048 24080 10100 24132
rect 41236 24080 41288 24132
rect 43444 24148 43496 24200
rect 43812 24191 43864 24200
rect 43812 24157 43821 24191
rect 43821 24157 43855 24191
rect 43855 24157 43864 24191
rect 43812 24148 43864 24157
rect 44180 24080 44232 24132
rect 45376 24123 45428 24132
rect 45376 24089 45403 24123
rect 45403 24089 45428 24123
rect 45376 24080 45428 24089
rect 53012 24284 53064 24336
rect 51632 24216 51684 24268
rect 55772 24216 55824 24268
rect 46664 24148 46716 24200
rect 46848 24191 46900 24200
rect 46848 24157 46857 24191
rect 46857 24157 46891 24191
rect 46891 24157 46900 24191
rect 46848 24148 46900 24157
rect 50804 24191 50856 24200
rect 50804 24157 50813 24191
rect 50813 24157 50847 24191
rect 50847 24157 50856 24191
rect 50804 24148 50856 24157
rect 52736 24148 52788 24200
rect 53104 24148 53156 24200
rect 53932 24148 53984 24200
rect 54668 24191 54720 24200
rect 54668 24157 54677 24191
rect 54677 24157 54711 24191
rect 54711 24157 54720 24191
rect 54668 24148 54720 24157
rect 55496 24191 55548 24200
rect 55496 24157 55505 24191
rect 55505 24157 55539 24191
rect 55539 24157 55548 24191
rect 55496 24148 55548 24157
rect 46940 24080 46992 24132
rect 52552 24080 52604 24132
rect 54760 24080 54812 24132
rect 56416 24148 56468 24200
rect 56968 24191 57020 24200
rect 56968 24157 56977 24191
rect 56977 24157 57011 24191
rect 57011 24157 57020 24191
rect 56968 24148 57020 24157
rect 57888 24148 57940 24200
rect 58072 24191 58124 24200
rect 58072 24157 58081 24191
rect 58081 24157 58115 24191
rect 58115 24157 58124 24191
rect 58072 24148 58124 24157
rect 56876 24080 56928 24132
rect 27804 24012 27856 24064
rect 39212 24012 39264 24064
rect 40224 24012 40276 24064
rect 44824 24012 44876 24064
rect 46848 24055 46900 24064
rect 46848 24021 46857 24055
rect 46857 24021 46891 24055
rect 46891 24021 46900 24055
rect 46848 24012 46900 24021
rect 56324 24012 56376 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 28724 23808 28776 23860
rect 31576 23851 31628 23860
rect 31576 23817 31585 23851
rect 31585 23817 31619 23851
rect 31619 23817 31628 23851
rect 31576 23808 31628 23817
rect 35256 23808 35308 23860
rect 36360 23851 36412 23860
rect 36360 23817 36369 23851
rect 36369 23817 36403 23851
rect 36403 23817 36412 23851
rect 36360 23808 36412 23817
rect 38752 23851 38804 23860
rect 38752 23817 38761 23851
rect 38761 23817 38795 23851
rect 38795 23817 38804 23851
rect 38752 23808 38804 23817
rect 39948 23851 40000 23860
rect 39948 23817 39957 23851
rect 39957 23817 39991 23851
rect 39991 23817 40000 23851
rect 39948 23808 40000 23817
rect 40224 23808 40276 23860
rect 30564 23740 30616 23792
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 25044 23672 25096 23724
rect 27528 23672 27580 23724
rect 27804 23715 27856 23724
rect 27804 23681 27813 23715
rect 27813 23681 27847 23715
rect 27847 23681 27856 23715
rect 27804 23672 27856 23681
rect 27988 23715 28040 23724
rect 27988 23681 27997 23715
rect 27997 23681 28031 23715
rect 28031 23681 28040 23715
rect 27988 23672 28040 23681
rect 30196 23715 30248 23724
rect 30196 23681 30205 23715
rect 30205 23681 30239 23715
rect 30239 23681 30248 23715
rect 30196 23672 30248 23681
rect 36452 23740 36504 23792
rect 38476 23740 38528 23792
rect 35900 23715 35952 23724
rect 24400 23604 24452 23656
rect 31300 23604 31352 23656
rect 35900 23681 35909 23715
rect 35909 23681 35943 23715
rect 35943 23681 35952 23715
rect 35900 23672 35952 23681
rect 39120 23715 39172 23724
rect 34520 23604 34572 23656
rect 39120 23681 39129 23715
rect 39129 23681 39163 23715
rect 39163 23681 39172 23715
rect 39120 23672 39172 23681
rect 40224 23715 40276 23724
rect 40224 23681 40234 23715
rect 40234 23681 40268 23715
rect 40268 23681 40276 23715
rect 40224 23672 40276 23681
rect 40592 23672 40644 23724
rect 40132 23647 40184 23656
rect 40132 23613 40141 23647
rect 40141 23613 40175 23647
rect 40175 23613 40184 23647
rect 40132 23604 40184 23613
rect 41236 23672 41288 23724
rect 42892 23808 42944 23860
rect 43904 23808 43956 23860
rect 43444 23740 43496 23792
rect 44180 23672 44232 23724
rect 44456 23715 44508 23724
rect 44456 23681 44465 23715
rect 44465 23681 44499 23715
rect 44499 23681 44508 23715
rect 44456 23672 44508 23681
rect 46020 23808 46072 23860
rect 46848 23808 46900 23860
rect 49884 23851 49936 23860
rect 46204 23740 46256 23792
rect 48596 23783 48648 23792
rect 48596 23749 48605 23783
rect 48605 23749 48639 23783
rect 48639 23749 48648 23783
rect 48596 23740 48648 23749
rect 48964 23740 49016 23792
rect 49884 23817 49893 23851
rect 49893 23817 49927 23851
rect 49927 23817 49936 23851
rect 49884 23808 49936 23817
rect 50804 23851 50856 23860
rect 50804 23817 50813 23851
rect 50813 23817 50847 23851
rect 50847 23817 50856 23851
rect 50804 23808 50856 23817
rect 53104 23851 53156 23860
rect 53104 23817 53113 23851
rect 53113 23817 53147 23851
rect 53147 23817 53156 23851
rect 53104 23808 53156 23817
rect 54208 23851 54260 23860
rect 54208 23817 54217 23851
rect 54217 23817 54251 23851
rect 54251 23817 54260 23851
rect 54208 23808 54260 23817
rect 56416 23851 56468 23860
rect 56416 23817 56425 23851
rect 56425 23817 56459 23851
rect 56459 23817 56468 23851
rect 56416 23808 56468 23817
rect 58164 23851 58216 23860
rect 58164 23817 58173 23851
rect 58173 23817 58207 23851
rect 58207 23817 58216 23851
rect 58164 23808 58216 23817
rect 50068 23740 50120 23792
rect 46664 23715 46716 23724
rect 46664 23681 46673 23715
rect 46673 23681 46707 23715
rect 46707 23681 46716 23715
rect 46664 23672 46716 23681
rect 46756 23715 46808 23724
rect 46756 23681 46765 23715
rect 46765 23681 46799 23715
rect 46799 23681 46808 23715
rect 46940 23715 46992 23724
rect 46756 23672 46808 23681
rect 46940 23681 46949 23715
rect 46949 23681 46983 23715
rect 46983 23681 46992 23715
rect 46940 23672 46992 23681
rect 47308 23672 47360 23724
rect 49700 23715 49752 23724
rect 49700 23681 49709 23715
rect 49709 23681 49743 23715
rect 49743 23681 49752 23715
rect 49700 23672 49752 23681
rect 49976 23672 50028 23724
rect 52000 23740 52052 23792
rect 51632 23672 51684 23724
rect 52092 23715 52144 23724
rect 52092 23681 52101 23715
rect 52101 23681 52135 23715
rect 52135 23681 52144 23715
rect 52092 23672 52144 23681
rect 52184 23715 52236 23724
rect 52184 23681 52193 23715
rect 52193 23681 52227 23715
rect 52227 23681 52236 23715
rect 53012 23715 53064 23724
rect 52184 23672 52236 23681
rect 53012 23681 53021 23715
rect 53021 23681 53055 23715
rect 53055 23681 53064 23715
rect 53012 23672 53064 23681
rect 53288 23672 53340 23724
rect 53840 23715 53892 23724
rect 53840 23681 53849 23715
rect 53849 23681 53883 23715
rect 53883 23681 53892 23715
rect 53840 23672 53892 23681
rect 56324 23715 56376 23724
rect 56324 23681 56333 23715
rect 56333 23681 56367 23715
rect 56367 23681 56376 23715
rect 56324 23672 56376 23681
rect 56416 23672 56468 23724
rect 48596 23604 48648 23656
rect 49424 23647 49476 23656
rect 49424 23613 49433 23647
rect 49433 23613 49467 23647
rect 49467 23613 49476 23647
rect 49424 23604 49476 23613
rect 53932 23647 53984 23656
rect 53932 23613 53941 23647
rect 53941 23613 53975 23647
rect 53975 23613 53984 23647
rect 53932 23604 53984 23613
rect 58164 23672 58216 23724
rect 57428 23604 57480 23656
rect 56876 23536 56928 23588
rect 1676 23511 1728 23520
rect 1676 23477 1685 23511
rect 1685 23477 1719 23511
rect 1719 23477 1728 23511
rect 1676 23468 1728 23477
rect 40868 23468 40920 23520
rect 41696 23511 41748 23520
rect 41696 23477 41705 23511
rect 41705 23477 41739 23511
rect 41739 23477 41748 23511
rect 41696 23468 41748 23477
rect 41972 23468 42024 23520
rect 44456 23468 44508 23520
rect 48688 23468 48740 23520
rect 49240 23468 49292 23520
rect 49792 23468 49844 23520
rect 51908 23468 51960 23520
rect 52460 23468 52512 23520
rect 57796 23468 57848 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 27528 23264 27580 23316
rect 30196 23264 30248 23316
rect 34520 23264 34572 23316
rect 35900 23264 35952 23316
rect 38476 23264 38528 23316
rect 39120 23264 39172 23316
rect 43444 23307 43496 23316
rect 43444 23273 43453 23307
rect 43453 23273 43487 23307
rect 43487 23273 43496 23307
rect 43444 23264 43496 23273
rect 45744 23264 45796 23316
rect 46664 23264 46716 23316
rect 49148 23264 49200 23316
rect 50160 23264 50212 23316
rect 52092 23307 52144 23316
rect 52092 23273 52101 23307
rect 52101 23273 52135 23307
rect 52135 23273 52144 23307
rect 52092 23264 52144 23273
rect 53196 23264 53248 23316
rect 53288 23264 53340 23316
rect 53840 23264 53892 23316
rect 57612 23307 57664 23316
rect 57612 23273 57621 23307
rect 57621 23273 57655 23307
rect 57655 23273 57664 23307
rect 57612 23264 57664 23273
rect 58072 23264 58124 23316
rect 28632 23239 28684 23248
rect 28632 23205 28641 23239
rect 28641 23205 28675 23239
rect 28675 23205 28684 23239
rect 28632 23196 28684 23205
rect 31024 23196 31076 23248
rect 22836 23060 22888 23112
rect 23388 23060 23440 23112
rect 32496 23128 32548 23180
rect 36452 23128 36504 23180
rect 45008 23196 45060 23248
rect 45560 23196 45612 23248
rect 49700 23239 49752 23248
rect 49700 23205 49709 23239
rect 49709 23205 49743 23239
rect 49743 23205 49752 23239
rect 49700 23196 49752 23205
rect 49976 23196 50028 23248
rect 56140 23196 56192 23248
rect 26240 23060 26292 23112
rect 26700 23103 26752 23112
rect 26700 23069 26709 23103
rect 26709 23069 26743 23103
rect 26743 23069 26752 23103
rect 26700 23060 26752 23069
rect 27068 23103 27120 23112
rect 27068 23069 27077 23103
rect 27077 23069 27111 23103
rect 27111 23069 27120 23103
rect 27068 23060 27120 23069
rect 27528 23060 27580 23112
rect 27988 23103 28040 23112
rect 27988 23069 27997 23103
rect 27997 23069 28031 23103
rect 28031 23069 28040 23103
rect 27988 23060 28040 23069
rect 29000 23060 29052 23112
rect 30564 23060 30616 23112
rect 30748 23103 30800 23112
rect 30748 23069 30757 23103
rect 30757 23069 30791 23103
rect 30791 23069 30800 23103
rect 30748 23060 30800 23069
rect 31668 23103 31720 23112
rect 31668 23069 31677 23103
rect 31677 23069 31711 23103
rect 31711 23069 31720 23103
rect 31668 23060 31720 23069
rect 28540 22992 28592 23044
rect 29460 22992 29512 23044
rect 32128 23060 32180 23112
rect 35348 23060 35400 23112
rect 36268 23103 36320 23112
rect 36268 23069 36277 23103
rect 36277 23069 36311 23103
rect 36311 23069 36320 23103
rect 36268 23060 36320 23069
rect 37464 23128 37516 23180
rect 41972 23171 42024 23180
rect 37280 23103 37332 23112
rect 37280 23069 37289 23103
rect 37289 23069 37323 23103
rect 37323 23069 37332 23103
rect 37280 23060 37332 23069
rect 38108 23103 38160 23112
rect 38108 23069 38117 23103
rect 38117 23069 38151 23103
rect 38151 23069 38160 23103
rect 38108 23060 38160 23069
rect 38292 23060 38344 23112
rect 41972 23137 41981 23171
rect 41981 23137 42015 23171
rect 42015 23137 42024 23171
rect 41972 23128 42024 23137
rect 44364 23171 44416 23180
rect 44364 23137 44373 23171
rect 44373 23137 44407 23171
rect 44407 23137 44416 23171
rect 44364 23128 44416 23137
rect 40500 23103 40552 23112
rect 34704 22992 34756 23044
rect 36728 22992 36780 23044
rect 40500 23069 40509 23103
rect 40509 23069 40543 23103
rect 40543 23069 40552 23103
rect 40500 23060 40552 23069
rect 40868 23103 40920 23112
rect 40868 23069 40877 23103
rect 40877 23069 40911 23103
rect 40911 23069 40920 23103
rect 40868 23060 40920 23069
rect 41604 23060 41656 23112
rect 44272 23103 44324 23112
rect 44272 23069 44281 23103
rect 44281 23069 44315 23103
rect 44315 23069 44324 23103
rect 44272 23060 44324 23069
rect 44640 23060 44692 23112
rect 45560 23103 45612 23112
rect 45560 23069 45569 23103
rect 45569 23069 45603 23103
rect 45603 23069 45612 23103
rect 45560 23060 45612 23069
rect 46020 23060 46072 23112
rect 15936 22924 15988 22976
rect 30288 22924 30340 22976
rect 31852 22924 31904 22976
rect 33968 22924 34020 22976
rect 38108 22924 38160 22976
rect 42432 22992 42484 23044
rect 48044 23128 48096 23180
rect 55588 23171 55640 23180
rect 46756 23060 46808 23112
rect 55588 23137 55597 23171
rect 55597 23137 55631 23171
rect 55631 23137 55640 23171
rect 55588 23128 55640 23137
rect 48688 23103 48740 23112
rect 48688 23069 48697 23103
rect 48697 23069 48731 23103
rect 48731 23069 48740 23103
rect 48688 23060 48740 23069
rect 48964 23103 49016 23112
rect 48964 23069 48973 23103
rect 48973 23069 49007 23103
rect 49007 23069 49016 23103
rect 48964 23060 49016 23069
rect 49792 23103 49844 23112
rect 49792 23069 49801 23103
rect 49801 23069 49835 23103
rect 49835 23069 49844 23103
rect 49792 23060 49844 23069
rect 49424 22992 49476 23044
rect 52184 23060 52236 23112
rect 55680 23103 55732 23112
rect 55680 23069 55689 23103
rect 55689 23069 55723 23103
rect 55723 23069 55732 23103
rect 55680 23060 55732 23069
rect 58256 23103 58308 23112
rect 44548 22924 44600 22976
rect 48596 22924 48648 22976
rect 53012 22992 53064 23044
rect 53196 22992 53248 23044
rect 54668 22992 54720 23044
rect 56968 22992 57020 23044
rect 57428 23035 57480 23044
rect 57428 23001 57437 23035
rect 57437 23001 57471 23035
rect 57471 23001 57480 23035
rect 58256 23069 58265 23103
rect 58265 23069 58299 23103
rect 58299 23069 58308 23103
rect 58256 23060 58308 23069
rect 57428 22992 57480 23001
rect 52000 22924 52052 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 27068 22720 27120 22772
rect 29000 22763 29052 22772
rect 29000 22729 29009 22763
rect 29009 22729 29043 22763
rect 29043 22729 29052 22763
rect 29000 22720 29052 22729
rect 37740 22720 37792 22772
rect 40500 22763 40552 22772
rect 2412 22652 2464 22704
rect 37280 22652 37332 22704
rect 39028 22652 39080 22704
rect 40500 22729 40509 22763
rect 40509 22729 40543 22763
rect 40543 22729 40552 22763
rect 40500 22720 40552 22729
rect 41696 22720 41748 22772
rect 42432 22720 42484 22772
rect 42892 22695 42944 22704
rect 26700 22584 26752 22636
rect 28816 22627 28868 22636
rect 28816 22593 28825 22627
rect 28825 22593 28859 22627
rect 28859 22593 28868 22627
rect 29460 22627 29512 22636
rect 28816 22584 28868 22593
rect 29460 22593 29469 22627
rect 29469 22593 29503 22627
rect 29503 22593 29512 22627
rect 29460 22584 29512 22593
rect 22836 22516 22888 22568
rect 26240 22516 26292 22568
rect 26976 22516 27028 22568
rect 27528 22516 27580 22568
rect 28540 22559 28592 22568
rect 28540 22525 28549 22559
rect 28549 22525 28583 22559
rect 28583 22525 28592 22559
rect 28540 22516 28592 22525
rect 23388 22448 23440 22500
rect 25044 22448 25096 22500
rect 23112 22423 23164 22432
rect 23112 22389 23121 22423
rect 23121 22389 23155 22423
rect 23155 22389 23164 22423
rect 23112 22380 23164 22389
rect 25872 22380 25924 22432
rect 30288 22627 30340 22636
rect 30288 22593 30297 22627
rect 30297 22593 30331 22627
rect 30331 22593 30340 22627
rect 30288 22584 30340 22593
rect 30564 22584 30616 22636
rect 31024 22627 31076 22636
rect 31024 22593 31033 22627
rect 31033 22593 31067 22627
rect 31067 22593 31076 22627
rect 31024 22584 31076 22593
rect 31300 22627 31352 22636
rect 31300 22593 31309 22627
rect 31309 22593 31343 22627
rect 31343 22593 31352 22627
rect 31300 22584 31352 22593
rect 31852 22584 31904 22636
rect 33968 22627 34020 22636
rect 33968 22593 33977 22627
rect 33977 22593 34011 22627
rect 34011 22593 34020 22627
rect 33968 22584 34020 22593
rect 34796 22627 34848 22636
rect 34796 22593 34805 22627
rect 34805 22593 34839 22627
rect 34839 22593 34848 22627
rect 34796 22584 34848 22593
rect 37464 22627 37516 22636
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 39212 22584 39264 22636
rect 39120 22448 39172 22500
rect 40132 22584 40184 22636
rect 40500 22627 40552 22636
rect 40500 22593 40509 22627
rect 40509 22593 40543 22627
rect 40543 22593 40552 22627
rect 40500 22584 40552 22593
rect 42892 22661 42901 22695
rect 42901 22661 42935 22695
rect 42935 22661 42944 22695
rect 42892 22652 42944 22661
rect 44180 22720 44232 22772
rect 46020 22720 46072 22772
rect 46664 22720 46716 22772
rect 48044 22763 48096 22772
rect 48044 22729 48053 22763
rect 48053 22729 48087 22763
rect 48087 22729 48096 22763
rect 48044 22720 48096 22729
rect 52000 22720 52052 22772
rect 56968 22763 57020 22772
rect 56968 22729 56977 22763
rect 56977 22729 57011 22763
rect 57011 22729 57020 22763
rect 56968 22720 57020 22729
rect 58164 22763 58216 22772
rect 58164 22729 58173 22763
rect 58173 22729 58207 22763
rect 58207 22729 58216 22763
rect 58164 22720 58216 22729
rect 46756 22652 46808 22704
rect 47308 22652 47360 22704
rect 40776 22584 40828 22636
rect 41328 22627 41380 22636
rect 41328 22593 41337 22627
rect 41337 22593 41371 22627
rect 41371 22593 41380 22627
rect 41328 22584 41380 22593
rect 45744 22627 45796 22636
rect 45744 22593 45753 22627
rect 45753 22593 45787 22627
rect 45787 22593 45796 22627
rect 45744 22584 45796 22593
rect 46204 22584 46256 22636
rect 46572 22584 46624 22636
rect 49240 22584 49292 22636
rect 51264 22584 51316 22636
rect 51724 22627 51776 22636
rect 51724 22593 51733 22627
rect 51733 22593 51767 22627
rect 51767 22593 51776 22627
rect 51724 22584 51776 22593
rect 53380 22627 53432 22636
rect 53380 22593 53389 22627
rect 53389 22593 53423 22627
rect 53423 22593 53432 22627
rect 53380 22584 53432 22593
rect 53564 22627 53616 22636
rect 53564 22593 53573 22627
rect 53573 22593 53607 22627
rect 53607 22593 53616 22627
rect 53564 22584 53616 22593
rect 53748 22584 53800 22636
rect 54668 22652 54720 22704
rect 56600 22695 56652 22704
rect 56600 22661 56609 22695
rect 56609 22661 56643 22695
rect 56643 22661 56652 22695
rect 56600 22652 56652 22661
rect 56784 22695 56836 22704
rect 56784 22661 56809 22695
rect 56809 22661 56836 22695
rect 56784 22652 56836 22661
rect 55128 22627 55180 22636
rect 40592 22516 40644 22568
rect 41604 22516 41656 22568
rect 45652 22559 45704 22568
rect 41512 22380 41564 22432
rect 45652 22525 45661 22559
rect 45661 22525 45695 22559
rect 45695 22525 45704 22559
rect 45652 22516 45704 22525
rect 45560 22448 45612 22500
rect 46112 22559 46164 22568
rect 46112 22525 46121 22559
rect 46121 22525 46155 22559
rect 46155 22525 46164 22559
rect 46112 22516 46164 22525
rect 49700 22516 49752 22568
rect 52092 22559 52144 22568
rect 52092 22525 52101 22559
rect 52101 22525 52135 22559
rect 52135 22525 52144 22559
rect 52092 22516 52144 22525
rect 52184 22516 52236 22568
rect 53656 22516 53708 22568
rect 55128 22593 55137 22627
rect 55137 22593 55171 22627
rect 55171 22593 55180 22627
rect 55128 22584 55180 22593
rect 55588 22627 55640 22636
rect 55588 22593 55597 22627
rect 55597 22593 55631 22627
rect 55631 22593 55640 22627
rect 55588 22584 55640 22593
rect 55864 22516 55916 22568
rect 52644 22448 52696 22500
rect 47676 22380 47728 22432
rect 49424 22380 49476 22432
rect 55680 22423 55732 22432
rect 55680 22389 55689 22423
rect 55689 22389 55723 22423
rect 55723 22389 55732 22423
rect 55680 22380 55732 22389
rect 56508 22380 56560 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 27528 22219 27580 22228
rect 27528 22185 27537 22219
rect 27537 22185 27571 22219
rect 27571 22185 27580 22219
rect 27528 22176 27580 22185
rect 23112 21972 23164 22024
rect 23388 21972 23440 22024
rect 24768 22040 24820 22092
rect 25044 22083 25096 22092
rect 25044 22049 25053 22083
rect 25053 22049 25087 22083
rect 25087 22049 25096 22083
rect 25044 22040 25096 22049
rect 28632 22176 28684 22228
rect 30748 22219 30800 22228
rect 30748 22185 30757 22219
rect 30757 22185 30791 22219
rect 30791 22185 30800 22219
rect 30748 22176 30800 22185
rect 34796 22176 34848 22228
rect 42432 22176 42484 22228
rect 44364 22176 44416 22228
rect 44548 22176 44600 22228
rect 32588 22108 32640 22160
rect 23756 21947 23808 21956
rect 23756 21913 23765 21947
rect 23765 21913 23799 21947
rect 23799 21913 23808 21947
rect 23756 21904 23808 21913
rect 24032 22015 24084 22024
rect 24032 21981 24041 22015
rect 24041 21981 24075 22015
rect 24075 21981 24084 22015
rect 24032 21972 24084 21981
rect 24676 21972 24728 22024
rect 25688 21972 25740 22024
rect 25872 21972 25924 22024
rect 26424 21972 26476 22024
rect 27068 22015 27120 22024
rect 27068 21981 27077 22015
rect 27077 21981 27111 22015
rect 27111 21981 27120 22015
rect 27068 21972 27120 21981
rect 27160 22015 27212 22024
rect 27160 21981 27169 22015
rect 27169 21981 27203 22015
rect 27203 21981 27212 22015
rect 27160 21972 27212 21981
rect 27712 21972 27764 22024
rect 31116 22015 31168 22024
rect 31116 21981 31125 22015
rect 31125 21981 31159 22015
rect 31159 21981 31168 22015
rect 31116 21972 31168 21981
rect 31300 21972 31352 22024
rect 31852 22040 31904 22092
rect 31760 22015 31812 22024
rect 31760 21981 31769 22015
rect 31769 21981 31803 22015
rect 31803 21981 31812 22015
rect 34520 22040 34572 22092
rect 38936 22040 38988 22092
rect 31760 21972 31812 21981
rect 32128 22015 32180 22024
rect 32128 21981 32137 22015
rect 32137 21981 32171 22015
rect 32171 21981 32180 22015
rect 32128 21972 32180 21981
rect 33324 21972 33376 22024
rect 35532 22015 35584 22024
rect 35532 21981 35541 22015
rect 35541 21981 35575 22015
rect 35575 21981 35584 22015
rect 35532 21972 35584 21981
rect 39028 22015 39080 22024
rect 31944 21947 31996 21956
rect 31944 21913 31953 21947
rect 31953 21913 31987 21947
rect 31987 21913 31996 21947
rect 31944 21904 31996 21913
rect 35440 21904 35492 21956
rect 39028 21981 39037 22015
rect 39037 21981 39071 22015
rect 39071 21981 39080 22015
rect 39028 21972 39080 21981
rect 39304 22015 39356 22024
rect 39304 21981 39313 22015
rect 39313 21981 39347 22015
rect 39347 21981 39356 22015
rect 39304 21972 39356 21981
rect 40500 22040 40552 22092
rect 40776 22040 40828 22092
rect 40960 22040 41012 22092
rect 45560 22108 45612 22160
rect 46296 22108 46348 22160
rect 48964 22176 49016 22228
rect 53104 22176 53156 22228
rect 53288 22219 53340 22228
rect 53288 22185 53297 22219
rect 53297 22185 53331 22219
rect 53331 22185 53340 22219
rect 53288 22176 53340 22185
rect 57428 22176 57480 22228
rect 58072 22176 58124 22228
rect 57980 22108 58032 22160
rect 41144 22015 41196 22024
rect 41144 21981 41153 22015
rect 41153 21981 41187 22015
rect 41187 21981 41196 22015
rect 47768 22040 47820 22092
rect 47860 22040 47912 22092
rect 49240 22083 49292 22092
rect 49240 22049 49249 22083
rect 49249 22049 49283 22083
rect 49283 22049 49292 22083
rect 49240 22040 49292 22049
rect 49424 22040 49476 22092
rect 50160 22040 50212 22092
rect 53564 22083 53616 22092
rect 53564 22049 53573 22083
rect 53573 22049 53607 22083
rect 53607 22049 53616 22083
rect 53564 22040 53616 22049
rect 55864 22083 55916 22092
rect 55864 22049 55873 22083
rect 55873 22049 55907 22083
rect 55907 22049 55916 22083
rect 55864 22040 55916 22049
rect 57796 22083 57848 22092
rect 57796 22049 57805 22083
rect 57805 22049 57839 22083
rect 57839 22049 57848 22083
rect 57796 22040 57848 22049
rect 41696 22015 41748 22024
rect 41144 21972 41196 21981
rect 41696 21981 41705 22015
rect 41705 21981 41739 22015
rect 41739 21981 41748 22015
rect 41696 21972 41748 21981
rect 40776 21947 40828 21956
rect 23848 21879 23900 21888
rect 23848 21845 23863 21879
rect 23863 21845 23897 21879
rect 23897 21845 23900 21879
rect 23848 21836 23900 21845
rect 24492 21836 24544 21888
rect 24860 21836 24912 21888
rect 26056 21836 26108 21888
rect 26240 21879 26292 21888
rect 26240 21845 26249 21879
rect 26249 21845 26283 21879
rect 26283 21845 26292 21879
rect 26240 21836 26292 21845
rect 31760 21836 31812 21888
rect 38936 21836 38988 21888
rect 39120 21879 39172 21888
rect 39120 21845 39129 21879
rect 39129 21845 39163 21879
rect 39163 21845 39172 21879
rect 39120 21836 39172 21845
rect 40224 21836 40276 21888
rect 40776 21913 40785 21947
rect 40785 21913 40819 21947
rect 40819 21913 40828 21947
rect 40776 21904 40828 21913
rect 40868 21947 40920 21956
rect 40868 21913 40877 21947
rect 40877 21913 40911 21947
rect 40911 21913 40920 21947
rect 40868 21904 40920 21913
rect 41328 21904 41380 21956
rect 40684 21836 40736 21888
rect 44824 21972 44876 22024
rect 45744 21972 45796 22024
rect 47124 22015 47176 22024
rect 47124 21981 47133 22015
rect 47133 21981 47167 22015
rect 47167 21981 47176 22015
rect 47124 21972 47176 21981
rect 48780 21972 48832 22024
rect 49148 22015 49200 22024
rect 49148 21981 49157 22015
rect 49157 21981 49191 22015
rect 49191 21981 49200 22015
rect 49148 21972 49200 21981
rect 50068 21972 50120 22024
rect 53380 21972 53432 22024
rect 53656 22015 53708 22024
rect 53656 21981 53665 22015
rect 53665 21981 53699 22015
rect 53699 21981 53708 22015
rect 53656 21972 53708 21981
rect 53748 22015 53800 22024
rect 53748 21981 53757 22015
rect 53757 21981 53791 22015
rect 53791 21981 53800 22015
rect 53748 21972 53800 21981
rect 44456 21947 44508 21956
rect 44456 21913 44465 21947
rect 44465 21913 44499 21947
rect 44499 21913 44508 21947
rect 44456 21904 44508 21913
rect 52644 21947 52696 21956
rect 52644 21913 52653 21947
rect 52653 21913 52687 21947
rect 52687 21913 52696 21947
rect 52644 21904 52696 21913
rect 52828 21947 52880 21956
rect 52828 21913 52837 21947
rect 52837 21913 52871 21947
rect 52871 21913 52880 21947
rect 52828 21904 52880 21913
rect 53104 21904 53156 21956
rect 54392 21904 54444 21956
rect 42156 21879 42208 21888
rect 42156 21845 42165 21879
rect 42165 21845 42199 21879
rect 42199 21845 42208 21879
rect 42156 21836 42208 21845
rect 44916 21836 44968 21888
rect 45376 21836 45428 21888
rect 46572 21836 46624 21888
rect 54300 21836 54352 21888
rect 55220 21972 55272 22024
rect 56508 22015 56560 22024
rect 56508 21981 56517 22015
rect 56517 21981 56551 22015
rect 56551 21981 56560 22015
rect 56508 21972 56560 21981
rect 58164 21972 58216 22024
rect 55036 21904 55088 21956
rect 56784 21947 56836 21956
rect 56784 21913 56793 21947
rect 56793 21913 56827 21947
rect 56827 21913 56836 21947
rect 56784 21904 56836 21913
rect 55128 21836 55180 21888
rect 56600 21879 56652 21888
rect 56600 21845 56609 21879
rect 56609 21845 56643 21879
rect 56643 21845 56652 21879
rect 56600 21836 56652 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 24492 21675 24544 21684
rect 24492 21641 24501 21675
rect 24501 21641 24535 21675
rect 24535 21641 24544 21675
rect 24492 21632 24544 21641
rect 24860 21675 24912 21684
rect 24860 21641 24869 21675
rect 24869 21641 24903 21675
rect 24903 21641 24912 21675
rect 24860 21632 24912 21641
rect 26240 21632 26292 21684
rect 27160 21632 27212 21684
rect 27712 21675 27764 21684
rect 27712 21641 27721 21675
rect 27721 21641 27755 21675
rect 27755 21641 27764 21675
rect 27712 21632 27764 21641
rect 31668 21632 31720 21684
rect 32128 21632 32180 21684
rect 36728 21632 36780 21684
rect 39304 21632 39356 21684
rect 40868 21632 40920 21684
rect 41236 21675 41288 21684
rect 41236 21641 41245 21675
rect 41245 21641 41279 21675
rect 41279 21641 41288 21675
rect 41236 21632 41288 21641
rect 47768 21675 47820 21684
rect 47768 21641 47777 21675
rect 47777 21641 47811 21675
rect 47811 21641 47820 21675
rect 47768 21632 47820 21641
rect 48780 21675 48832 21684
rect 48780 21641 48789 21675
rect 48789 21641 48823 21675
rect 48823 21641 48832 21675
rect 48780 21632 48832 21641
rect 49240 21632 49292 21684
rect 50068 21632 50120 21684
rect 52828 21632 52880 21684
rect 54392 21632 54444 21684
rect 55128 21675 55180 21684
rect 55128 21641 55137 21675
rect 55137 21641 55171 21675
rect 55171 21641 55180 21675
rect 55128 21632 55180 21641
rect 56784 21632 56836 21684
rect 58164 21675 58216 21684
rect 58164 21641 58173 21675
rect 58173 21641 58207 21675
rect 58207 21641 58216 21675
rect 58164 21632 58216 21641
rect 24032 21564 24084 21616
rect 23664 21496 23716 21548
rect 23756 21496 23808 21548
rect 24768 21496 24820 21548
rect 24952 21539 25004 21548
rect 24952 21505 24961 21539
rect 24961 21505 24995 21539
rect 24995 21505 25004 21539
rect 24952 21496 25004 21505
rect 25044 21496 25096 21548
rect 27436 21564 27488 21616
rect 30564 21607 30616 21616
rect 30564 21573 30573 21607
rect 30573 21573 30607 21607
rect 30607 21573 30616 21607
rect 30564 21564 30616 21573
rect 31944 21564 31996 21616
rect 26056 21496 26108 21548
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 28080 21539 28132 21548
rect 28080 21505 28089 21539
rect 28089 21505 28123 21539
rect 28123 21505 28132 21539
rect 28080 21496 28132 21505
rect 30012 21539 30064 21548
rect 30012 21505 30021 21539
rect 30021 21505 30055 21539
rect 30055 21505 30064 21539
rect 30012 21496 30064 21505
rect 30472 21539 30524 21548
rect 30472 21505 30481 21539
rect 30481 21505 30515 21539
rect 30515 21505 30524 21539
rect 30472 21496 30524 21505
rect 30656 21539 30708 21548
rect 30656 21505 30665 21539
rect 30665 21505 30699 21539
rect 30699 21505 30708 21539
rect 30656 21496 30708 21505
rect 31116 21496 31168 21548
rect 22192 21428 22244 21480
rect 23388 21471 23440 21480
rect 23388 21437 23397 21471
rect 23397 21437 23431 21471
rect 23431 21437 23440 21471
rect 23388 21428 23440 21437
rect 27712 21428 27764 21480
rect 31300 21428 31352 21480
rect 31760 21539 31812 21548
rect 31760 21505 31769 21539
rect 31769 21505 31803 21539
rect 31803 21505 31812 21539
rect 31760 21496 31812 21505
rect 32220 21496 32272 21548
rect 33692 21539 33744 21548
rect 33692 21505 33701 21539
rect 33701 21505 33735 21539
rect 33735 21505 33744 21539
rect 33692 21496 33744 21505
rect 35440 21564 35492 21616
rect 35532 21539 35584 21548
rect 32588 21471 32640 21480
rect 32588 21437 32597 21471
rect 32597 21437 32631 21471
rect 32631 21437 32640 21471
rect 32588 21428 32640 21437
rect 32956 21428 33008 21480
rect 35532 21505 35541 21539
rect 35541 21505 35575 21539
rect 35575 21505 35584 21539
rect 35532 21496 35584 21505
rect 35900 21496 35952 21548
rect 36636 21539 36688 21548
rect 36636 21505 36645 21539
rect 36645 21505 36679 21539
rect 36679 21505 36688 21539
rect 36636 21496 36688 21505
rect 37372 21496 37424 21548
rect 37556 21471 37608 21480
rect 37556 21437 37565 21471
rect 37565 21437 37599 21471
rect 37599 21437 37608 21471
rect 37556 21428 37608 21437
rect 38200 21496 38252 21548
rect 40684 21564 40736 21616
rect 42064 21564 42116 21616
rect 42156 21564 42208 21616
rect 43720 21607 43772 21616
rect 40592 21496 40644 21548
rect 38476 21428 38528 21480
rect 41052 21428 41104 21480
rect 43720 21573 43729 21607
rect 43729 21573 43763 21607
rect 43763 21573 43772 21607
rect 43720 21564 43772 21573
rect 44456 21564 44508 21616
rect 45284 21564 45336 21616
rect 46572 21564 46624 21616
rect 47768 21539 47820 21548
rect 47768 21505 47777 21539
rect 47777 21505 47811 21539
rect 47811 21505 47820 21539
rect 47768 21496 47820 21505
rect 47860 21496 47912 21548
rect 48228 21496 48280 21548
rect 49240 21496 49292 21548
rect 54484 21564 54536 21616
rect 54392 21539 54444 21548
rect 54392 21505 54401 21539
rect 54401 21505 54435 21539
rect 54435 21505 54444 21539
rect 54392 21496 54444 21505
rect 55036 21539 55088 21548
rect 55036 21505 55045 21539
rect 55045 21505 55079 21539
rect 55079 21505 55088 21539
rect 55036 21496 55088 21505
rect 55220 21539 55272 21548
rect 55220 21505 55229 21539
rect 55229 21505 55263 21539
rect 55263 21505 55272 21539
rect 55220 21496 55272 21505
rect 56876 21539 56928 21548
rect 56876 21505 56885 21539
rect 56885 21505 56919 21539
rect 56919 21505 56928 21539
rect 56876 21496 56928 21505
rect 56968 21496 57020 21548
rect 57888 21496 57940 21548
rect 58348 21496 58400 21548
rect 43444 21428 43496 21480
rect 25504 21335 25556 21344
rect 25504 21301 25513 21335
rect 25513 21301 25547 21335
rect 25547 21301 25556 21335
rect 25504 21292 25556 21301
rect 25688 21292 25740 21344
rect 32312 21360 32364 21412
rect 28632 21292 28684 21344
rect 32956 21292 33008 21344
rect 33784 21335 33836 21344
rect 33784 21301 33793 21335
rect 33793 21301 33827 21335
rect 33827 21301 33836 21335
rect 33784 21292 33836 21301
rect 43168 21292 43220 21344
rect 46940 21335 46992 21344
rect 46940 21301 46949 21335
rect 46949 21301 46983 21335
rect 46983 21301 46992 21335
rect 46940 21292 46992 21301
rect 48964 21335 49016 21344
rect 48964 21301 48973 21335
rect 48973 21301 49007 21335
rect 49007 21301 49016 21335
rect 48964 21292 49016 21301
rect 54576 21292 54628 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 23664 21131 23716 21140
rect 23664 21097 23673 21131
rect 23673 21097 23707 21131
rect 23707 21097 23716 21131
rect 23664 21088 23716 21097
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 23848 20884 23900 20893
rect 24676 21088 24728 21140
rect 24952 21088 25004 21140
rect 27896 21088 27948 21140
rect 28080 21088 28132 21140
rect 30288 21088 30340 21140
rect 31484 21131 31536 21140
rect 31484 21097 31493 21131
rect 31493 21097 31527 21131
rect 31527 21097 31536 21131
rect 31484 21088 31536 21097
rect 32312 21131 32364 21140
rect 32312 21097 32321 21131
rect 32321 21097 32355 21131
rect 32355 21097 32364 21131
rect 32312 21088 32364 21097
rect 33324 21131 33376 21140
rect 33324 21097 33333 21131
rect 33333 21097 33367 21131
rect 33367 21097 33376 21131
rect 33324 21088 33376 21097
rect 35900 21131 35952 21140
rect 35900 21097 35909 21131
rect 35909 21097 35943 21131
rect 35943 21097 35952 21131
rect 35900 21088 35952 21097
rect 38108 21088 38160 21140
rect 38292 21088 38344 21140
rect 45744 21088 45796 21140
rect 46940 21088 46992 21140
rect 49148 21088 49200 21140
rect 54392 21088 54444 21140
rect 56876 21131 56928 21140
rect 56876 21097 56885 21131
rect 56885 21097 56919 21131
rect 56919 21097 56928 21131
rect 56876 21088 56928 21097
rect 56968 21088 57020 21140
rect 57888 21131 57940 21140
rect 57888 21097 57897 21131
rect 57897 21097 57931 21131
rect 57931 21097 57940 21131
rect 57888 21088 57940 21097
rect 26056 20952 26108 21004
rect 27712 20952 27764 21004
rect 26148 20927 26200 20936
rect 26148 20893 26157 20927
rect 26157 20893 26191 20927
rect 26191 20893 26200 20927
rect 26148 20884 26200 20893
rect 24768 20859 24820 20868
rect 24768 20825 24795 20859
rect 24795 20825 24820 20859
rect 24768 20816 24820 20825
rect 24860 20816 24912 20868
rect 25504 20816 25556 20868
rect 26424 20927 26476 20936
rect 26424 20893 26433 20927
rect 26433 20893 26467 20927
rect 26467 20893 26476 20927
rect 28448 20927 28500 20936
rect 26424 20884 26476 20893
rect 28448 20893 28457 20927
rect 28457 20893 28491 20927
rect 28491 20893 28500 20927
rect 28448 20884 28500 20893
rect 28540 20816 28592 20868
rect 27804 20791 27856 20800
rect 27804 20757 27829 20791
rect 27829 20757 27856 20791
rect 30012 20927 30064 20936
rect 30012 20893 30021 20927
rect 30021 20893 30055 20927
rect 30055 20893 30064 20927
rect 30012 20884 30064 20893
rect 30656 20952 30708 21004
rect 30932 20952 30984 21004
rect 30472 20884 30524 20936
rect 31300 20884 31352 20936
rect 30564 20816 30616 20868
rect 31576 20884 31628 20936
rect 33692 21020 33744 21072
rect 35532 21020 35584 21072
rect 42432 21020 42484 21072
rect 47492 21063 47544 21072
rect 47492 21029 47501 21063
rect 47501 21029 47535 21063
rect 47535 21029 47544 21063
rect 47492 21020 47544 21029
rect 52552 21063 52604 21072
rect 52552 21029 52561 21063
rect 52561 21029 52595 21063
rect 52595 21029 52604 21063
rect 52552 21020 52604 21029
rect 33784 20952 33836 21004
rect 35716 20952 35768 21004
rect 38200 20995 38252 21004
rect 38200 20961 38209 20995
rect 38209 20961 38243 20995
rect 38243 20961 38252 20995
rect 38200 20952 38252 20961
rect 43260 20952 43312 21004
rect 51264 20952 51316 21004
rect 52000 20952 52052 21004
rect 34520 20884 34572 20936
rect 35532 20927 35584 20936
rect 35532 20893 35541 20927
rect 35541 20893 35575 20927
rect 35575 20893 35584 20927
rect 35532 20884 35584 20893
rect 37372 20927 37424 20936
rect 32956 20859 33008 20868
rect 32956 20825 32965 20859
rect 32965 20825 32999 20859
rect 32999 20825 33008 20859
rect 32956 20816 33008 20825
rect 33508 20816 33560 20868
rect 37372 20893 37381 20927
rect 37381 20893 37415 20927
rect 37415 20893 37424 20927
rect 37372 20884 37424 20893
rect 37556 20927 37608 20936
rect 37556 20893 37565 20927
rect 37565 20893 37599 20927
rect 37599 20893 37608 20927
rect 37556 20884 37608 20893
rect 38476 20884 38528 20936
rect 42432 20884 42484 20936
rect 47952 20927 48004 20936
rect 43168 20859 43220 20868
rect 27804 20748 27856 20757
rect 32220 20748 32272 20800
rect 35624 20748 35676 20800
rect 36636 20748 36688 20800
rect 39396 20748 39448 20800
rect 42616 20748 42668 20800
rect 43168 20825 43177 20859
rect 43177 20825 43211 20859
rect 43211 20825 43220 20859
rect 43168 20816 43220 20825
rect 47952 20893 47961 20927
rect 47961 20893 47995 20927
rect 47995 20893 48004 20927
rect 47952 20884 48004 20893
rect 48136 20927 48188 20936
rect 48136 20893 48145 20927
rect 48145 20893 48179 20927
rect 48179 20893 48188 20927
rect 48136 20884 48188 20893
rect 48228 20884 48280 20936
rect 48964 20884 49016 20936
rect 49148 20927 49200 20936
rect 49148 20893 49157 20927
rect 49157 20893 49191 20927
rect 49191 20893 49200 20927
rect 49148 20884 49200 20893
rect 50896 20884 50948 20936
rect 51356 20927 51408 20936
rect 51356 20893 51365 20927
rect 51365 20893 51399 20927
rect 51399 20893 51408 20927
rect 51356 20884 51408 20893
rect 51540 20927 51592 20936
rect 51540 20893 51549 20927
rect 51549 20893 51583 20927
rect 51583 20893 51592 20927
rect 51540 20884 51592 20893
rect 53012 20927 53064 20936
rect 53012 20893 53021 20927
rect 53021 20893 53055 20927
rect 53055 20893 53064 20927
rect 53012 20884 53064 20893
rect 53288 20927 53340 20936
rect 53288 20893 53297 20927
rect 53297 20893 53331 20927
rect 53331 20893 53340 20927
rect 53288 20884 53340 20893
rect 47400 20816 47452 20868
rect 44548 20748 44600 20800
rect 45284 20748 45336 20800
rect 45744 20748 45796 20800
rect 55496 21020 55548 21072
rect 55404 20952 55456 21004
rect 53840 20884 53892 20936
rect 54024 20884 54076 20936
rect 54300 20927 54352 20936
rect 54300 20893 54309 20927
rect 54309 20893 54343 20927
rect 54343 20893 54352 20927
rect 54300 20884 54352 20893
rect 54576 20884 54628 20936
rect 55680 20884 55732 20936
rect 56508 20859 56560 20868
rect 56508 20825 56517 20859
rect 56517 20825 56551 20859
rect 56551 20825 56560 20859
rect 56508 20816 56560 20825
rect 57520 20859 57572 20868
rect 56600 20748 56652 20800
rect 57520 20825 57529 20859
rect 57529 20825 57563 20859
rect 57563 20825 57572 20859
rect 57520 20816 57572 20825
rect 57704 20791 57756 20800
rect 57704 20757 57729 20791
rect 57729 20757 57756 20791
rect 57704 20748 57756 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 24768 20544 24820 20596
rect 25688 20587 25740 20596
rect 25688 20553 25697 20587
rect 25697 20553 25731 20587
rect 25731 20553 25740 20587
rect 25688 20544 25740 20553
rect 26240 20587 26292 20596
rect 26240 20553 26249 20587
rect 26249 20553 26283 20587
rect 26283 20553 26292 20587
rect 26240 20544 26292 20553
rect 26332 20544 26384 20596
rect 28448 20544 28500 20596
rect 28540 20544 28592 20596
rect 30472 20587 30524 20596
rect 30472 20553 30481 20587
rect 30481 20553 30515 20587
rect 30515 20553 30524 20587
rect 30472 20544 30524 20553
rect 31484 20587 31536 20596
rect 31484 20553 31493 20587
rect 31493 20553 31527 20587
rect 31527 20553 31536 20587
rect 31484 20544 31536 20553
rect 22836 20519 22888 20528
rect 22836 20485 22845 20519
rect 22845 20485 22879 20519
rect 22879 20485 22888 20519
rect 22836 20476 22888 20485
rect 23296 20476 23348 20528
rect 28632 20519 28684 20528
rect 28632 20485 28641 20519
rect 28641 20485 28675 20519
rect 28675 20485 28684 20519
rect 28632 20476 28684 20485
rect 23572 20451 23624 20460
rect 23572 20417 23581 20451
rect 23581 20417 23615 20451
rect 23615 20417 23624 20451
rect 23572 20408 23624 20417
rect 24032 20408 24084 20460
rect 25504 20451 25556 20460
rect 25504 20417 25513 20451
rect 25513 20417 25547 20451
rect 25547 20417 25556 20451
rect 25504 20408 25556 20417
rect 26424 20408 26476 20460
rect 26608 20451 26660 20460
rect 26608 20417 26617 20451
rect 26617 20417 26651 20451
rect 26651 20417 26660 20451
rect 27896 20451 27948 20460
rect 26608 20408 26660 20417
rect 27896 20417 27905 20451
rect 27905 20417 27939 20451
rect 27939 20417 27948 20451
rect 27896 20408 27948 20417
rect 29736 20408 29788 20460
rect 30564 20408 30616 20460
rect 31300 20476 31352 20528
rect 33692 20544 33744 20596
rect 34520 20544 34572 20596
rect 41052 20587 41104 20596
rect 30932 20451 30984 20460
rect 30932 20417 30941 20451
rect 30941 20417 30975 20451
rect 30975 20417 30984 20451
rect 30932 20408 30984 20417
rect 31392 20451 31444 20460
rect 31392 20417 31401 20451
rect 31401 20417 31435 20451
rect 31435 20417 31444 20451
rect 31392 20408 31444 20417
rect 31668 20451 31720 20460
rect 31668 20417 31677 20451
rect 31677 20417 31711 20451
rect 31711 20417 31720 20451
rect 31668 20408 31720 20417
rect 31760 20451 31812 20460
rect 31760 20417 31769 20451
rect 31769 20417 31803 20451
rect 31803 20417 31812 20451
rect 31760 20408 31812 20417
rect 33232 20408 33284 20460
rect 33416 20451 33468 20460
rect 33416 20417 33425 20451
rect 33425 20417 33459 20451
rect 33459 20417 33468 20451
rect 33416 20408 33468 20417
rect 33784 20408 33836 20460
rect 35440 20451 35492 20460
rect 35440 20417 35449 20451
rect 35449 20417 35483 20451
rect 35483 20417 35492 20451
rect 35440 20408 35492 20417
rect 36728 20408 36780 20460
rect 36912 20408 36964 20460
rect 38844 20451 38896 20460
rect 38844 20417 38853 20451
rect 38853 20417 38887 20451
rect 38887 20417 38896 20451
rect 38844 20408 38896 20417
rect 41052 20553 41061 20587
rect 41061 20553 41095 20587
rect 41095 20553 41104 20587
rect 41052 20544 41104 20553
rect 43444 20544 43496 20596
rect 48964 20544 49016 20596
rect 47952 20476 48004 20528
rect 53288 20544 53340 20596
rect 40040 20408 40092 20460
rect 41236 20408 41288 20460
rect 41696 20451 41748 20460
rect 41696 20417 41705 20451
rect 41705 20417 41739 20451
rect 41739 20417 41748 20451
rect 41696 20408 41748 20417
rect 41880 20408 41932 20460
rect 42616 20451 42668 20460
rect 42616 20417 42625 20451
rect 42625 20417 42659 20451
rect 42659 20417 42668 20451
rect 42616 20408 42668 20417
rect 44456 20451 44508 20460
rect 44456 20417 44465 20451
rect 44465 20417 44499 20451
rect 44499 20417 44508 20451
rect 44456 20408 44508 20417
rect 24492 20383 24544 20392
rect 24492 20349 24501 20383
rect 24501 20349 24535 20383
rect 24535 20349 24544 20383
rect 24492 20340 24544 20349
rect 23940 20272 23992 20324
rect 29276 20340 29328 20392
rect 31484 20340 31536 20392
rect 26516 20272 26568 20324
rect 27528 20272 27580 20324
rect 32220 20340 32272 20392
rect 35992 20340 36044 20392
rect 38752 20383 38804 20392
rect 38752 20349 38761 20383
rect 38761 20349 38795 20383
rect 38795 20349 38804 20383
rect 38752 20340 38804 20349
rect 40316 20383 40368 20392
rect 40316 20349 40325 20383
rect 40325 20349 40359 20383
rect 40359 20349 40368 20383
rect 40316 20340 40368 20349
rect 44364 20383 44416 20392
rect 44364 20349 44373 20383
rect 44373 20349 44407 20383
rect 44407 20349 44416 20383
rect 44364 20340 44416 20349
rect 45560 20408 45612 20460
rect 48136 20408 48188 20460
rect 48780 20408 48832 20460
rect 49792 20476 49844 20528
rect 50896 20476 50948 20528
rect 50068 20451 50120 20460
rect 45744 20340 45796 20392
rect 50068 20417 50077 20451
rect 50077 20417 50111 20451
rect 50111 20417 50120 20451
rect 50068 20408 50120 20417
rect 50160 20451 50212 20460
rect 50160 20417 50169 20451
rect 50169 20417 50203 20451
rect 50203 20417 50212 20451
rect 51080 20476 51132 20528
rect 51540 20476 51592 20528
rect 55220 20544 55272 20596
rect 57520 20544 57572 20596
rect 54760 20519 54812 20528
rect 54760 20485 54769 20519
rect 54769 20485 54803 20519
rect 54803 20485 54812 20519
rect 54760 20476 54812 20485
rect 56968 20476 57020 20528
rect 57704 20476 57756 20528
rect 50160 20408 50212 20417
rect 51172 20451 51224 20460
rect 51172 20417 51181 20451
rect 51181 20417 51215 20451
rect 51215 20417 51224 20451
rect 51172 20408 51224 20417
rect 48872 20272 48924 20324
rect 50896 20340 50948 20392
rect 52552 20408 52604 20460
rect 52736 20340 52788 20392
rect 54024 20408 54076 20460
rect 54208 20408 54260 20460
rect 53196 20383 53248 20392
rect 53196 20349 53205 20383
rect 53205 20349 53239 20383
rect 53239 20349 53248 20383
rect 53196 20340 53248 20349
rect 54484 20451 54536 20460
rect 54484 20417 54510 20451
rect 54510 20417 54536 20451
rect 54484 20408 54536 20417
rect 55404 20408 55456 20460
rect 56600 20451 56652 20460
rect 56600 20417 56609 20451
rect 56609 20417 56643 20451
rect 56643 20417 56652 20451
rect 56600 20408 56652 20417
rect 56508 20340 56560 20392
rect 54484 20272 54536 20324
rect 58348 20315 58400 20324
rect 58348 20281 58357 20315
rect 58357 20281 58391 20315
rect 58391 20281 58400 20315
rect 58348 20272 58400 20281
rect 36084 20247 36136 20256
rect 36084 20213 36093 20247
rect 36093 20213 36127 20247
rect 36127 20213 36136 20247
rect 36084 20204 36136 20213
rect 36728 20204 36780 20256
rect 41420 20204 41472 20256
rect 42800 20247 42852 20256
rect 42800 20213 42809 20247
rect 42809 20213 42843 20247
rect 42843 20213 42852 20247
rect 42800 20204 42852 20213
rect 49148 20247 49200 20256
rect 49148 20213 49157 20247
rect 49157 20213 49191 20247
rect 49191 20213 49200 20247
rect 49148 20204 49200 20213
rect 51816 20204 51868 20256
rect 53012 20247 53064 20256
rect 53012 20213 53021 20247
rect 53021 20213 53055 20247
rect 53055 20213 53064 20247
rect 53012 20204 53064 20213
rect 54300 20204 54352 20256
rect 54760 20204 54812 20256
rect 55680 20247 55732 20256
rect 55680 20213 55689 20247
rect 55689 20213 55723 20247
rect 55723 20213 55732 20247
rect 55680 20204 55732 20213
rect 56692 20204 56744 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 23572 20000 23624 20052
rect 23940 20043 23992 20052
rect 23940 20009 23949 20043
rect 23949 20009 23983 20043
rect 23983 20009 23992 20043
rect 23940 20000 23992 20009
rect 27068 20043 27120 20052
rect 27068 20009 27077 20043
rect 27077 20009 27111 20043
rect 27111 20009 27120 20043
rect 27068 20000 27120 20009
rect 28264 20000 28316 20052
rect 29736 20043 29788 20052
rect 26516 19975 26568 19984
rect 26516 19941 26525 19975
rect 26525 19941 26559 19975
rect 26559 19941 26568 19975
rect 26516 19932 26568 19941
rect 27988 19932 28040 19984
rect 24492 19864 24544 19916
rect 25504 19907 25556 19916
rect 25504 19873 25513 19907
rect 25513 19873 25547 19907
rect 25547 19873 25556 19907
rect 25504 19864 25556 19873
rect 28264 19907 28316 19916
rect 24032 19839 24084 19848
rect 24032 19805 24041 19839
rect 24041 19805 24075 19839
rect 24075 19805 24084 19839
rect 24032 19796 24084 19805
rect 25320 19839 25372 19848
rect 25320 19805 25329 19839
rect 25329 19805 25363 19839
rect 25363 19805 25372 19839
rect 25320 19796 25372 19805
rect 26240 19796 26292 19848
rect 26424 19796 26476 19848
rect 28264 19873 28273 19907
rect 28273 19873 28307 19907
rect 28307 19873 28316 19907
rect 28264 19864 28316 19873
rect 28632 19932 28684 19984
rect 29736 20009 29745 20043
rect 29745 20009 29779 20043
rect 29779 20009 29788 20043
rect 29736 20000 29788 20009
rect 31668 20000 31720 20052
rect 33508 20043 33560 20052
rect 33508 20009 33517 20043
rect 33517 20009 33551 20043
rect 33551 20009 33560 20043
rect 33508 20000 33560 20009
rect 35440 20000 35492 20052
rect 38844 20043 38896 20052
rect 38844 20009 38853 20043
rect 38853 20009 38887 20043
rect 38887 20009 38896 20043
rect 38844 20000 38896 20009
rect 39028 20000 39080 20052
rect 40592 20000 40644 20052
rect 44364 20043 44416 20052
rect 44364 20009 44373 20043
rect 44373 20009 44407 20043
rect 44407 20009 44416 20043
rect 44364 20000 44416 20009
rect 47124 20000 47176 20052
rect 47400 20043 47452 20052
rect 47400 20009 47409 20043
rect 47409 20009 47443 20043
rect 47443 20009 47452 20043
rect 47400 20000 47452 20009
rect 49148 20043 49200 20052
rect 49148 20009 49157 20043
rect 49157 20009 49191 20043
rect 49191 20009 49200 20043
rect 49148 20000 49200 20009
rect 51172 20000 51224 20052
rect 54208 20000 54260 20052
rect 56324 20000 56376 20052
rect 57704 20000 57756 20052
rect 38752 19932 38804 19984
rect 46296 19932 46348 19984
rect 47768 19975 47820 19984
rect 47768 19941 47777 19975
rect 47777 19941 47811 19975
rect 47811 19941 47820 19975
rect 47768 19932 47820 19941
rect 48596 19932 48648 19984
rect 54024 19932 54076 19984
rect 29276 19864 29328 19916
rect 28356 19839 28408 19848
rect 28356 19805 28365 19839
rect 28365 19805 28399 19839
rect 28399 19805 28408 19839
rect 28356 19796 28408 19805
rect 29920 19839 29972 19848
rect 25044 19728 25096 19780
rect 26608 19728 26660 19780
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 29552 19728 29604 19780
rect 31576 19796 31628 19848
rect 32220 19796 32272 19848
rect 33416 19864 33468 19916
rect 36544 19907 36596 19916
rect 34612 19796 34664 19848
rect 35808 19796 35860 19848
rect 36544 19873 36553 19907
rect 36553 19873 36587 19907
rect 36587 19873 36596 19907
rect 36544 19864 36596 19873
rect 36728 19907 36780 19916
rect 36728 19873 36737 19907
rect 36737 19873 36771 19907
rect 36771 19873 36780 19907
rect 36728 19864 36780 19873
rect 38016 19864 38068 19916
rect 37464 19796 37516 19848
rect 37832 19839 37884 19848
rect 37832 19805 37841 19839
rect 37841 19805 37875 19839
rect 37875 19805 37884 19839
rect 37832 19796 37884 19805
rect 40040 19907 40092 19916
rect 40040 19873 40049 19907
rect 40049 19873 40083 19907
rect 40083 19873 40092 19907
rect 40040 19864 40092 19873
rect 41420 19907 41472 19916
rect 41420 19873 41429 19907
rect 41429 19873 41463 19907
rect 41463 19873 41472 19907
rect 42800 19907 42852 19916
rect 41420 19864 41472 19873
rect 42800 19873 42809 19907
rect 42809 19873 42843 19907
rect 42843 19873 42852 19907
rect 42800 19864 42852 19873
rect 46020 19864 46072 19916
rect 40316 19796 40368 19848
rect 41512 19796 41564 19848
rect 43076 19839 43128 19848
rect 43076 19805 43085 19839
rect 43085 19805 43119 19839
rect 43119 19805 43128 19839
rect 43076 19796 43128 19805
rect 33232 19728 33284 19780
rect 33784 19728 33836 19780
rect 36084 19728 36136 19780
rect 42248 19771 42300 19780
rect 42248 19737 42257 19771
rect 42257 19737 42291 19771
rect 42291 19737 42300 19771
rect 42248 19728 42300 19737
rect 26332 19660 26384 19712
rect 28080 19703 28132 19712
rect 28080 19669 28089 19703
rect 28089 19669 28123 19703
rect 28123 19669 28132 19703
rect 28080 19660 28132 19669
rect 28540 19660 28592 19712
rect 30932 19660 30984 19712
rect 32680 19660 32732 19712
rect 36820 19703 36872 19712
rect 36820 19669 36829 19703
rect 36829 19669 36863 19703
rect 36863 19669 36872 19703
rect 36820 19660 36872 19669
rect 43720 19660 43772 19712
rect 44548 19796 44600 19848
rect 45560 19839 45612 19848
rect 45560 19805 45569 19839
rect 45569 19805 45603 19839
rect 45603 19805 45612 19839
rect 45560 19796 45612 19805
rect 45744 19839 45796 19848
rect 45744 19805 45753 19839
rect 45753 19805 45787 19839
rect 45787 19805 45796 19839
rect 45744 19796 45796 19805
rect 45652 19728 45704 19780
rect 48964 19864 49016 19916
rect 52828 19864 52880 19916
rect 47492 19728 47544 19780
rect 48228 19796 48280 19848
rect 48872 19839 48924 19848
rect 48872 19805 48881 19839
rect 48881 19805 48915 19839
rect 48915 19805 48924 19839
rect 48872 19796 48924 19805
rect 48596 19728 48648 19780
rect 50896 19796 50948 19848
rect 49148 19728 49200 19780
rect 51080 19839 51132 19848
rect 51080 19805 51089 19839
rect 51089 19805 51123 19839
rect 51123 19805 51132 19839
rect 52000 19839 52052 19848
rect 51080 19796 51132 19805
rect 52000 19805 52009 19839
rect 52009 19805 52043 19839
rect 52043 19805 52052 19839
rect 52000 19796 52052 19805
rect 52736 19796 52788 19848
rect 53104 19796 53156 19848
rect 53564 19864 53616 19916
rect 54760 19864 54812 19916
rect 56600 19907 56652 19916
rect 56600 19873 56609 19907
rect 56609 19873 56643 19907
rect 56643 19873 56652 19907
rect 56600 19864 56652 19873
rect 57428 19907 57480 19916
rect 57428 19873 57437 19907
rect 57437 19873 57471 19907
rect 57471 19873 57480 19907
rect 57428 19864 57480 19873
rect 54116 19839 54168 19848
rect 53288 19728 53340 19780
rect 54116 19805 54125 19839
rect 54125 19805 54159 19839
rect 54159 19805 54168 19839
rect 54116 19796 54168 19805
rect 54300 19796 54352 19848
rect 54484 19839 54536 19848
rect 54484 19805 54493 19839
rect 54493 19805 54527 19839
rect 54527 19805 54536 19839
rect 54484 19796 54536 19805
rect 55496 19839 55548 19848
rect 55496 19805 55505 19839
rect 55505 19805 55539 19839
rect 55539 19805 55548 19839
rect 55496 19796 55548 19805
rect 55404 19728 55456 19780
rect 56508 19796 56560 19848
rect 47860 19660 47912 19712
rect 51080 19660 51132 19712
rect 52092 19703 52144 19712
rect 52092 19669 52101 19703
rect 52101 19669 52135 19703
rect 52135 19669 52144 19703
rect 52092 19660 52144 19669
rect 53380 19660 53432 19712
rect 54024 19660 54076 19712
rect 55496 19660 55548 19712
rect 56416 19660 56468 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 23756 19499 23808 19508
rect 23756 19465 23765 19499
rect 23765 19465 23799 19499
rect 23799 19465 23808 19499
rect 23756 19456 23808 19465
rect 25044 19456 25096 19508
rect 25504 19499 25556 19508
rect 25504 19465 25513 19499
rect 25513 19465 25547 19499
rect 25547 19465 25556 19499
rect 25504 19456 25556 19465
rect 26056 19499 26108 19508
rect 26056 19465 26065 19499
rect 26065 19465 26099 19499
rect 26099 19465 26108 19499
rect 26056 19456 26108 19465
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 25412 19363 25464 19372
rect 23848 19252 23900 19304
rect 25412 19329 25421 19363
rect 25421 19329 25455 19363
rect 25455 19329 25464 19363
rect 25412 19320 25464 19329
rect 28632 19388 28684 19440
rect 34612 19456 34664 19508
rect 34704 19456 34756 19508
rect 36912 19499 36964 19508
rect 36912 19465 36921 19499
rect 36921 19465 36955 19499
rect 36955 19465 36964 19499
rect 36912 19456 36964 19465
rect 39120 19456 39172 19508
rect 41236 19499 41288 19508
rect 41236 19465 41245 19499
rect 41245 19465 41279 19499
rect 41279 19465 41288 19499
rect 41236 19456 41288 19465
rect 41880 19499 41932 19508
rect 41880 19465 41889 19499
rect 41889 19465 41923 19499
rect 41923 19465 41932 19499
rect 41880 19456 41932 19465
rect 43076 19456 43128 19508
rect 43720 19499 43772 19508
rect 43720 19465 43729 19499
rect 43729 19465 43763 19499
rect 43763 19465 43772 19499
rect 43720 19456 43772 19465
rect 48228 19456 48280 19508
rect 48596 19456 48648 19508
rect 28080 19363 28132 19372
rect 26240 19295 26292 19304
rect 26240 19261 26249 19295
rect 26249 19261 26283 19295
rect 26283 19261 26292 19295
rect 26240 19252 26292 19261
rect 26332 19295 26384 19304
rect 26332 19261 26341 19295
rect 26341 19261 26375 19295
rect 26375 19261 26384 19295
rect 26332 19252 26384 19261
rect 26516 19295 26568 19304
rect 26516 19261 26525 19295
rect 26525 19261 26559 19295
rect 26559 19261 26568 19295
rect 28080 19329 28089 19363
rect 28089 19329 28123 19363
rect 28123 19329 28132 19363
rect 28080 19320 28132 19329
rect 28356 19320 28408 19372
rect 28908 19363 28960 19372
rect 28908 19329 28917 19363
rect 28917 19329 28951 19363
rect 28951 19329 28960 19363
rect 28908 19320 28960 19329
rect 32680 19388 32732 19440
rect 29920 19363 29972 19372
rect 29920 19329 29929 19363
rect 29929 19329 29963 19363
rect 29963 19329 29972 19363
rect 29920 19320 29972 19329
rect 30380 19320 30432 19372
rect 31576 19363 31628 19372
rect 31576 19329 31585 19363
rect 31585 19329 31619 19363
rect 31619 19329 31628 19363
rect 31576 19320 31628 19329
rect 32220 19320 32272 19372
rect 32404 19320 32456 19372
rect 33140 19320 33192 19372
rect 34520 19388 34572 19440
rect 36360 19388 36412 19440
rect 39396 19431 39448 19440
rect 39396 19397 39405 19431
rect 39405 19397 39439 19431
rect 39439 19397 39448 19431
rect 39856 19431 39908 19440
rect 39396 19388 39448 19397
rect 39856 19397 39865 19431
rect 39865 19397 39899 19431
rect 39899 19397 39908 19431
rect 39856 19388 39908 19397
rect 40040 19431 40092 19440
rect 40040 19397 40065 19431
rect 40065 19397 40092 19431
rect 40040 19388 40092 19397
rect 45744 19388 45796 19440
rect 34428 19363 34480 19372
rect 34428 19329 34437 19363
rect 34437 19329 34471 19363
rect 34471 19329 34480 19363
rect 34428 19320 34480 19329
rect 26516 19252 26568 19261
rect 25136 19184 25188 19236
rect 27160 19252 27212 19304
rect 27712 19295 27764 19304
rect 27712 19261 27721 19295
rect 27721 19261 27755 19295
rect 27755 19261 27764 19295
rect 27712 19252 27764 19261
rect 29644 19252 29696 19304
rect 29828 19295 29880 19304
rect 29828 19261 29837 19295
rect 29837 19261 29871 19295
rect 29871 19261 29880 19295
rect 29828 19252 29880 19261
rect 29552 19184 29604 19236
rect 31852 19252 31904 19304
rect 32496 19295 32548 19304
rect 31760 19184 31812 19236
rect 32496 19261 32505 19295
rect 32505 19261 32539 19295
rect 32539 19261 32548 19295
rect 32496 19252 32548 19261
rect 33232 19252 33284 19304
rect 34888 19320 34940 19372
rect 35532 19363 35584 19372
rect 35532 19329 35541 19363
rect 35541 19329 35575 19363
rect 35575 19329 35584 19363
rect 35532 19320 35584 19329
rect 37832 19363 37884 19372
rect 34796 19252 34848 19304
rect 37832 19329 37841 19363
rect 37841 19329 37875 19363
rect 37875 19329 37884 19363
rect 37832 19320 37884 19329
rect 38016 19363 38068 19372
rect 38016 19329 38025 19363
rect 38025 19329 38059 19363
rect 38059 19329 38068 19363
rect 38016 19320 38068 19329
rect 41144 19363 41196 19372
rect 41144 19329 41153 19363
rect 41153 19329 41187 19363
rect 41187 19329 41196 19363
rect 41144 19320 41196 19329
rect 41420 19320 41472 19372
rect 41880 19320 41932 19372
rect 42800 19320 42852 19372
rect 43628 19363 43680 19372
rect 43628 19329 43637 19363
rect 43637 19329 43671 19363
rect 43671 19329 43680 19363
rect 43628 19320 43680 19329
rect 44088 19320 44140 19372
rect 46020 19363 46072 19372
rect 46020 19329 46029 19363
rect 46029 19329 46063 19363
rect 46063 19329 46072 19363
rect 46020 19320 46072 19329
rect 50160 19456 50212 19508
rect 51356 19499 51408 19508
rect 51356 19465 51365 19499
rect 51365 19465 51399 19499
rect 51399 19465 51408 19499
rect 51356 19456 51408 19465
rect 52092 19456 52144 19508
rect 53104 19499 53156 19508
rect 53104 19465 53113 19499
rect 53113 19465 53147 19499
rect 53147 19465 53156 19499
rect 53104 19456 53156 19465
rect 54944 19456 54996 19508
rect 57428 19456 57480 19508
rect 52000 19388 52052 19440
rect 43996 19252 44048 19304
rect 44548 19252 44600 19304
rect 45008 19295 45060 19304
rect 45008 19261 45017 19295
rect 45017 19261 45051 19295
rect 45051 19261 45060 19295
rect 45008 19252 45060 19261
rect 46296 19252 46348 19304
rect 46756 19252 46808 19304
rect 36544 19184 36596 19236
rect 36728 19227 36780 19236
rect 36728 19193 36737 19227
rect 36737 19193 36771 19227
rect 36771 19193 36780 19227
rect 36728 19184 36780 19193
rect 22100 19116 22152 19168
rect 25412 19116 25464 19168
rect 28540 19116 28592 19168
rect 40040 19159 40092 19168
rect 40040 19125 40049 19159
rect 40049 19125 40083 19159
rect 40083 19125 40092 19159
rect 40040 19116 40092 19125
rect 40224 19159 40276 19168
rect 40224 19125 40233 19159
rect 40233 19125 40267 19159
rect 40267 19125 40276 19159
rect 40224 19116 40276 19125
rect 43260 19159 43312 19168
rect 43260 19125 43269 19159
rect 43269 19125 43303 19159
rect 43303 19125 43312 19159
rect 43260 19116 43312 19125
rect 45836 19116 45888 19168
rect 50160 19363 50212 19372
rect 50160 19329 50169 19363
rect 50169 19329 50203 19363
rect 50203 19329 50212 19363
rect 50160 19320 50212 19329
rect 56048 19388 56100 19440
rect 53380 19363 53432 19372
rect 48136 19252 48188 19304
rect 49976 19295 50028 19304
rect 49976 19261 49985 19295
rect 49985 19261 50019 19295
rect 50019 19261 50028 19295
rect 49976 19252 50028 19261
rect 53380 19329 53389 19363
rect 53389 19329 53423 19363
rect 53423 19329 53432 19363
rect 53380 19320 53432 19329
rect 54116 19320 54168 19372
rect 56416 19320 56468 19372
rect 52000 19295 52052 19304
rect 48780 19184 48832 19236
rect 49148 19184 49200 19236
rect 52000 19261 52009 19295
rect 52009 19261 52043 19295
rect 52043 19261 52052 19295
rect 52000 19252 52052 19261
rect 53564 19252 53616 19304
rect 55496 19295 55548 19304
rect 55496 19261 55505 19295
rect 55505 19261 55539 19295
rect 55539 19261 55548 19295
rect 55496 19252 55548 19261
rect 55956 19252 56008 19304
rect 56600 19252 56652 19304
rect 50712 19116 50764 19168
rect 53288 19159 53340 19168
rect 53288 19125 53297 19159
rect 53297 19125 53331 19159
rect 53331 19125 53340 19159
rect 53288 19116 53340 19125
rect 53656 19116 53708 19168
rect 58348 19116 58400 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 22284 18912 22336 18964
rect 27528 18912 27580 18964
rect 29828 18912 29880 18964
rect 30564 18912 30616 18964
rect 31576 18955 31628 18964
rect 31576 18921 31585 18955
rect 31585 18921 31619 18955
rect 31619 18921 31628 18955
rect 31576 18912 31628 18921
rect 32496 18955 32548 18964
rect 32496 18921 32505 18955
rect 32505 18921 32539 18955
rect 32539 18921 32548 18955
rect 32496 18912 32548 18921
rect 34796 18912 34848 18964
rect 35624 18912 35676 18964
rect 37556 18912 37608 18964
rect 40040 18912 40092 18964
rect 40316 18912 40368 18964
rect 42800 18955 42852 18964
rect 42800 18921 42809 18955
rect 42809 18921 42843 18955
rect 42843 18921 42852 18955
rect 42800 18912 42852 18921
rect 46020 18912 46072 18964
rect 47492 18955 47544 18964
rect 47492 18921 47501 18955
rect 47501 18921 47535 18955
rect 47535 18921 47544 18955
rect 47492 18912 47544 18921
rect 51080 18955 51132 18964
rect 51080 18921 51089 18955
rect 51089 18921 51123 18955
rect 51123 18921 51132 18955
rect 55496 18955 55548 18964
rect 51080 18912 51132 18921
rect 55496 18921 55505 18955
rect 55505 18921 55539 18955
rect 55539 18921 55548 18955
rect 55496 18912 55548 18921
rect 26700 18844 26752 18896
rect 30012 18776 30064 18828
rect 23756 18708 23808 18760
rect 25136 18708 25188 18760
rect 25780 18708 25832 18760
rect 29276 18708 29328 18760
rect 30380 18751 30432 18760
rect 30380 18717 30389 18751
rect 30389 18717 30423 18751
rect 30423 18717 30432 18751
rect 30380 18708 30432 18717
rect 25688 18640 25740 18692
rect 26424 18683 26476 18692
rect 26424 18649 26433 18683
rect 26433 18649 26467 18683
rect 26467 18649 26476 18683
rect 26424 18640 26476 18649
rect 29092 18640 29144 18692
rect 32128 18708 32180 18760
rect 32220 18708 32272 18760
rect 32680 18751 32732 18760
rect 32680 18717 32689 18751
rect 32689 18717 32723 18751
rect 32723 18717 32732 18751
rect 32680 18708 32732 18717
rect 22284 18572 22336 18624
rect 23848 18572 23900 18624
rect 25596 18572 25648 18624
rect 33232 18776 33284 18828
rect 34520 18776 34572 18828
rect 35808 18819 35860 18828
rect 35808 18785 35817 18819
rect 35817 18785 35851 18819
rect 35851 18785 35860 18819
rect 35808 18776 35860 18785
rect 35992 18751 36044 18760
rect 35992 18717 36001 18751
rect 36001 18717 36035 18751
rect 36035 18717 36044 18751
rect 35992 18708 36044 18717
rect 36728 18751 36780 18760
rect 36728 18717 36737 18751
rect 36737 18717 36771 18751
rect 36771 18717 36780 18751
rect 36728 18708 36780 18717
rect 36912 18751 36964 18760
rect 36912 18717 36921 18751
rect 36921 18717 36955 18751
rect 36955 18717 36964 18751
rect 36912 18708 36964 18717
rect 35624 18640 35676 18692
rect 38660 18776 38712 18828
rect 39028 18844 39080 18896
rect 45008 18844 45060 18896
rect 39396 18776 39448 18828
rect 40132 18819 40184 18828
rect 40132 18785 40141 18819
rect 40141 18785 40175 18819
rect 40175 18785 40184 18819
rect 40132 18776 40184 18785
rect 40224 18776 40276 18828
rect 37832 18683 37884 18692
rect 37832 18649 37841 18683
rect 37841 18649 37875 18683
rect 37875 18649 37884 18683
rect 37832 18640 37884 18649
rect 39212 18708 39264 18760
rect 39304 18751 39356 18760
rect 39304 18717 39313 18751
rect 39313 18717 39347 18751
rect 39347 18717 39356 18751
rect 40592 18751 40644 18760
rect 39304 18708 39356 18717
rect 40592 18717 40601 18751
rect 40601 18717 40635 18751
rect 40635 18717 40644 18751
rect 40592 18708 40644 18717
rect 41788 18819 41840 18828
rect 36636 18572 36688 18624
rect 36728 18615 36780 18624
rect 36728 18581 36737 18615
rect 36737 18581 36771 18615
rect 36771 18581 36780 18615
rect 36728 18572 36780 18581
rect 37372 18572 37424 18624
rect 39580 18640 39632 18692
rect 41788 18785 41797 18819
rect 41797 18785 41831 18819
rect 41831 18785 41840 18819
rect 41788 18776 41840 18785
rect 45744 18776 45796 18828
rect 46388 18776 46440 18828
rect 49700 18776 49752 18828
rect 50988 18776 51040 18828
rect 51908 18844 51960 18896
rect 43260 18708 43312 18760
rect 46756 18708 46808 18760
rect 46940 18751 46992 18760
rect 46940 18717 46949 18751
rect 46949 18717 46983 18751
rect 46983 18717 46992 18751
rect 46940 18708 46992 18717
rect 47584 18751 47636 18760
rect 47584 18717 47593 18751
rect 47593 18717 47627 18751
rect 47627 18717 47636 18751
rect 47584 18708 47636 18717
rect 50160 18708 50212 18760
rect 50712 18751 50764 18760
rect 50712 18717 50721 18751
rect 50721 18717 50755 18751
rect 50755 18717 50764 18751
rect 50712 18708 50764 18717
rect 43168 18572 43220 18624
rect 52460 18708 52512 18760
rect 52920 18776 52972 18828
rect 55772 18819 55824 18828
rect 54024 18708 54076 18760
rect 43996 18572 44048 18624
rect 45744 18572 45796 18624
rect 45928 18615 45980 18624
rect 45928 18581 45937 18615
rect 45937 18581 45971 18615
rect 45971 18581 45980 18615
rect 45928 18572 45980 18581
rect 47216 18572 47268 18624
rect 50160 18572 50212 18624
rect 53932 18640 53984 18692
rect 55772 18785 55781 18819
rect 55781 18785 55815 18819
rect 55815 18785 55824 18819
rect 55772 18776 55824 18785
rect 55128 18708 55180 18760
rect 58348 18708 58400 18760
rect 55956 18640 56008 18692
rect 55680 18572 55732 18624
rect 56048 18572 56100 18624
rect 57244 18615 57296 18624
rect 57244 18581 57253 18615
rect 57253 18581 57287 18615
rect 57287 18581 57296 18615
rect 57244 18572 57296 18581
rect 58256 18615 58308 18624
rect 58256 18581 58265 18615
rect 58265 18581 58299 18615
rect 58299 18581 58308 18615
rect 58256 18572 58308 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 22100 18368 22152 18420
rect 23940 18368 23992 18420
rect 25044 18368 25096 18420
rect 26240 18368 26292 18420
rect 26332 18368 26384 18420
rect 27896 18368 27948 18420
rect 30012 18411 30064 18420
rect 30012 18377 30021 18411
rect 30021 18377 30055 18411
rect 30055 18377 30064 18411
rect 30012 18368 30064 18377
rect 31116 18368 31168 18420
rect 35256 18368 35308 18420
rect 35348 18368 35400 18420
rect 36728 18368 36780 18420
rect 38016 18368 38068 18420
rect 40132 18368 40184 18420
rect 41144 18368 41196 18420
rect 44272 18368 44324 18420
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 23848 18300 23900 18352
rect 24860 18343 24912 18352
rect 24860 18309 24869 18343
rect 24869 18309 24903 18343
rect 24903 18309 24912 18343
rect 24860 18300 24912 18309
rect 24768 18275 24820 18284
rect 24768 18241 24777 18275
rect 24777 18241 24811 18275
rect 24811 18241 24820 18275
rect 24768 18232 24820 18241
rect 22284 18207 22336 18216
rect 22284 18173 22293 18207
rect 22293 18173 22327 18207
rect 22327 18173 22336 18207
rect 22284 18164 22336 18173
rect 23296 18164 23348 18216
rect 25136 18232 25188 18284
rect 25504 18275 25556 18284
rect 25504 18241 25513 18275
rect 25513 18241 25547 18275
rect 25547 18241 25556 18275
rect 25504 18232 25556 18241
rect 25596 18275 25648 18284
rect 25596 18241 25605 18275
rect 25605 18241 25639 18275
rect 25639 18241 25648 18275
rect 26240 18275 26292 18284
rect 25596 18232 25648 18241
rect 26240 18241 26249 18275
rect 26249 18241 26283 18275
rect 26283 18241 26292 18275
rect 26240 18232 26292 18241
rect 26424 18300 26476 18352
rect 37372 18300 37424 18352
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 29552 18275 29604 18284
rect 29552 18241 29561 18275
rect 29561 18241 29595 18275
rect 29595 18241 29604 18275
rect 29552 18232 29604 18241
rect 29920 18232 29972 18284
rect 30472 18275 30524 18284
rect 30472 18241 30481 18275
rect 30481 18241 30515 18275
rect 30515 18241 30524 18275
rect 31116 18275 31168 18284
rect 30472 18232 30524 18241
rect 31116 18241 31125 18275
rect 31125 18241 31159 18275
rect 31159 18241 31168 18275
rect 31116 18232 31168 18241
rect 32772 18232 32824 18284
rect 32956 18275 33008 18284
rect 32956 18241 32965 18275
rect 32965 18241 32999 18275
rect 32999 18241 33008 18275
rect 33140 18275 33192 18284
rect 32956 18232 33008 18241
rect 33140 18241 33149 18275
rect 33149 18241 33183 18275
rect 33183 18241 33192 18275
rect 33140 18232 33192 18241
rect 27252 18164 27304 18216
rect 27896 18207 27948 18216
rect 27896 18173 27905 18207
rect 27905 18173 27939 18207
rect 27939 18173 27948 18207
rect 27896 18164 27948 18173
rect 28080 18207 28132 18216
rect 28080 18173 28089 18207
rect 28089 18173 28123 18207
rect 28123 18173 28132 18207
rect 28080 18164 28132 18173
rect 31852 18164 31904 18216
rect 32220 18164 32272 18216
rect 36544 18232 36596 18284
rect 36636 18232 36688 18284
rect 38384 18275 38436 18284
rect 38384 18241 38393 18275
rect 38393 18241 38427 18275
rect 38427 18241 38436 18275
rect 38384 18232 38436 18241
rect 39028 18232 39080 18284
rect 39580 18275 39632 18284
rect 39580 18241 39589 18275
rect 39589 18241 39623 18275
rect 39623 18241 39632 18275
rect 39580 18232 39632 18241
rect 41788 18300 41840 18352
rect 41420 18275 41472 18284
rect 41420 18241 41429 18275
rect 41429 18241 41463 18275
rect 41463 18241 41472 18275
rect 41420 18232 41472 18241
rect 43720 18232 43772 18284
rect 44456 18232 44508 18284
rect 45652 18275 45704 18284
rect 45652 18241 45661 18275
rect 45661 18241 45695 18275
rect 45695 18241 45704 18275
rect 45652 18232 45704 18241
rect 52184 18368 52236 18420
rect 52828 18368 52880 18420
rect 55128 18411 55180 18420
rect 55128 18377 55137 18411
rect 55137 18377 55171 18411
rect 55171 18377 55180 18411
rect 55128 18368 55180 18377
rect 46388 18343 46440 18352
rect 46388 18309 46397 18343
rect 46397 18309 46431 18343
rect 46431 18309 46440 18343
rect 46388 18300 46440 18309
rect 36728 18164 36780 18216
rect 37464 18207 37516 18216
rect 37464 18173 37473 18207
rect 37473 18173 37507 18207
rect 37507 18173 37516 18207
rect 37464 18164 37516 18173
rect 39212 18164 39264 18216
rect 44548 18164 44600 18216
rect 29644 18139 29696 18148
rect 1768 18071 1820 18080
rect 1768 18037 1777 18071
rect 1777 18037 1811 18071
rect 1811 18037 1820 18071
rect 1768 18028 1820 18037
rect 29644 18105 29653 18139
rect 29653 18105 29687 18139
rect 29687 18105 29696 18139
rect 29644 18096 29696 18105
rect 29828 18096 29880 18148
rect 44824 18164 44876 18216
rect 50712 18300 50764 18352
rect 53748 18343 53800 18352
rect 53748 18309 53757 18343
rect 53757 18309 53791 18343
rect 53791 18309 53800 18343
rect 53748 18300 53800 18309
rect 55680 18343 55732 18352
rect 55680 18309 55689 18343
rect 55689 18309 55723 18343
rect 55723 18309 55732 18343
rect 55680 18300 55732 18309
rect 48504 18275 48556 18284
rect 48504 18241 48513 18275
rect 48513 18241 48547 18275
rect 48547 18241 48556 18275
rect 48504 18232 48556 18241
rect 48964 18275 49016 18284
rect 48964 18241 48973 18275
rect 48973 18241 49007 18275
rect 49007 18241 49016 18275
rect 48964 18232 49016 18241
rect 50160 18275 50212 18284
rect 50160 18241 50169 18275
rect 50169 18241 50203 18275
rect 50203 18241 50212 18275
rect 50160 18232 50212 18241
rect 51908 18232 51960 18284
rect 27528 18028 27580 18080
rect 28264 18028 28316 18080
rect 28540 18028 28592 18080
rect 28908 18028 28960 18080
rect 35256 18028 35308 18080
rect 36912 18028 36964 18080
rect 37372 18028 37424 18080
rect 45008 18096 45060 18148
rect 51172 18164 51224 18216
rect 51448 18164 51500 18216
rect 53656 18275 53708 18284
rect 53656 18241 53665 18275
rect 53665 18241 53699 18275
rect 53699 18241 53708 18275
rect 53656 18232 53708 18241
rect 53932 18275 53984 18284
rect 53932 18241 53941 18275
rect 53941 18241 53975 18275
rect 53975 18241 53984 18275
rect 53932 18232 53984 18241
rect 55772 18275 55824 18284
rect 55772 18241 55781 18275
rect 55781 18241 55815 18275
rect 55815 18241 55824 18275
rect 55772 18232 55824 18241
rect 55956 18275 56008 18284
rect 55956 18241 55965 18275
rect 55965 18241 55999 18275
rect 55999 18241 56008 18275
rect 55956 18232 56008 18241
rect 57796 18232 57848 18284
rect 47584 18096 47636 18148
rect 49516 18096 49568 18148
rect 39304 18071 39356 18080
rect 39304 18037 39313 18071
rect 39313 18037 39347 18071
rect 39347 18037 39356 18071
rect 39304 18028 39356 18037
rect 43904 18071 43956 18080
rect 43904 18037 43913 18071
rect 43913 18037 43947 18071
rect 43947 18037 43956 18071
rect 43904 18028 43956 18037
rect 48412 18028 48464 18080
rect 49792 18028 49844 18080
rect 50160 18096 50212 18148
rect 50896 18139 50948 18148
rect 50896 18105 50905 18139
rect 50905 18105 50939 18139
rect 50939 18105 50948 18139
rect 50896 18096 50948 18105
rect 54208 18096 54260 18148
rect 57428 18096 57480 18148
rect 51908 18071 51960 18080
rect 51908 18037 51917 18071
rect 51917 18037 51951 18071
rect 51951 18037 51960 18071
rect 51908 18028 51960 18037
rect 52368 18028 52420 18080
rect 54760 18028 54812 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 23296 17867 23348 17876
rect 23296 17833 23305 17867
rect 23305 17833 23339 17867
rect 23339 17833 23348 17867
rect 23296 17824 23348 17833
rect 24032 17824 24084 17876
rect 24952 17824 25004 17876
rect 25780 17824 25832 17876
rect 27528 17824 27580 17876
rect 1584 17799 1636 17808
rect 1584 17765 1593 17799
rect 1593 17765 1627 17799
rect 1627 17765 1636 17799
rect 1584 17756 1636 17765
rect 27252 17756 27304 17808
rect 27804 17824 27856 17876
rect 33232 17824 33284 17876
rect 33784 17867 33836 17876
rect 33784 17833 33793 17867
rect 33793 17833 33827 17867
rect 33827 17833 33836 17867
rect 33784 17824 33836 17833
rect 35440 17824 35492 17876
rect 36452 17824 36504 17876
rect 24032 17731 24084 17740
rect 24032 17697 24041 17731
rect 24041 17697 24075 17731
rect 24075 17697 24084 17731
rect 24032 17688 24084 17697
rect 24768 17731 24820 17740
rect 24768 17697 24777 17731
rect 24777 17697 24811 17731
rect 24811 17697 24820 17731
rect 24768 17688 24820 17697
rect 24860 17731 24912 17740
rect 24860 17697 24869 17731
rect 24869 17697 24903 17731
rect 24903 17697 24912 17731
rect 24860 17688 24912 17697
rect 23756 17663 23808 17672
rect 23756 17629 23765 17663
rect 23765 17629 23799 17663
rect 23799 17629 23808 17663
rect 23756 17620 23808 17629
rect 25044 17663 25096 17672
rect 25044 17629 25053 17663
rect 25053 17629 25087 17663
rect 25087 17629 25096 17663
rect 25044 17620 25096 17629
rect 25136 17552 25188 17604
rect 25688 17552 25740 17604
rect 26240 17552 26292 17604
rect 26700 17620 26752 17672
rect 27528 17731 27580 17740
rect 27528 17697 27537 17731
rect 27537 17697 27571 17731
rect 27571 17697 27580 17731
rect 27528 17688 27580 17697
rect 31392 17756 31444 17808
rect 29092 17731 29144 17740
rect 29092 17697 29101 17731
rect 29101 17697 29135 17731
rect 29135 17697 29144 17731
rect 29092 17688 29144 17697
rect 31208 17688 31260 17740
rect 32312 17688 32364 17740
rect 34520 17756 34572 17808
rect 27988 17663 28040 17672
rect 27988 17629 27997 17663
rect 27997 17629 28031 17663
rect 28031 17629 28040 17663
rect 27988 17620 28040 17629
rect 28172 17620 28224 17672
rect 28264 17620 28316 17672
rect 30932 17663 30984 17672
rect 30932 17629 30941 17663
rect 30941 17629 30975 17663
rect 30975 17629 30984 17663
rect 30932 17620 30984 17629
rect 32404 17663 32456 17672
rect 32404 17629 32413 17663
rect 32413 17629 32447 17663
rect 32447 17629 32456 17663
rect 32404 17620 32456 17629
rect 32680 17620 32732 17672
rect 25596 17527 25648 17536
rect 25596 17493 25605 17527
rect 25605 17493 25639 17527
rect 25639 17493 25648 17527
rect 25596 17484 25648 17493
rect 32128 17552 32180 17604
rect 33232 17620 33284 17672
rect 34060 17688 34112 17740
rect 37740 17688 37792 17740
rect 33692 17663 33744 17672
rect 33692 17629 33701 17663
rect 33701 17629 33735 17663
rect 33735 17629 33744 17663
rect 33692 17620 33744 17629
rect 34520 17620 34572 17672
rect 36636 17620 36688 17672
rect 37188 17663 37240 17672
rect 37188 17629 37197 17663
rect 37197 17629 37231 17663
rect 37231 17629 37240 17663
rect 37188 17620 37240 17629
rect 37280 17663 37332 17672
rect 37280 17629 37289 17663
rect 37289 17629 37323 17663
rect 37323 17629 37332 17663
rect 37280 17620 37332 17629
rect 37464 17663 37516 17672
rect 37464 17629 37473 17663
rect 37473 17629 37507 17663
rect 37507 17629 37516 17663
rect 37464 17620 37516 17629
rect 38752 17824 38804 17876
rect 39212 17867 39264 17876
rect 39212 17833 39221 17867
rect 39221 17833 39255 17867
rect 39255 17833 39264 17867
rect 39212 17824 39264 17833
rect 44548 17824 44600 17876
rect 46020 17824 46072 17876
rect 44824 17756 44876 17808
rect 46112 17756 46164 17808
rect 47492 17824 47544 17876
rect 47768 17756 47820 17808
rect 48504 17824 48556 17876
rect 50988 17867 51040 17876
rect 50988 17833 50997 17867
rect 50997 17833 51031 17867
rect 51031 17833 51040 17867
rect 50988 17824 51040 17833
rect 51724 17824 51776 17876
rect 53104 17824 53156 17876
rect 53472 17824 53524 17876
rect 54484 17824 54536 17876
rect 55588 17824 55640 17876
rect 57796 17867 57848 17876
rect 57796 17833 57805 17867
rect 57805 17833 57839 17867
rect 57839 17833 57848 17867
rect 57796 17824 57848 17833
rect 48964 17756 49016 17808
rect 49792 17731 49844 17740
rect 43444 17663 43496 17672
rect 28080 17484 28132 17536
rect 28264 17484 28316 17536
rect 36636 17484 36688 17536
rect 38568 17552 38620 17604
rect 43444 17629 43453 17663
rect 43453 17629 43487 17663
rect 43487 17629 43496 17663
rect 43444 17620 43496 17629
rect 43536 17552 43588 17604
rect 43720 17663 43772 17672
rect 43720 17629 43729 17663
rect 43729 17629 43763 17663
rect 43763 17629 43772 17663
rect 43720 17620 43772 17629
rect 44180 17620 44232 17672
rect 45284 17620 45336 17672
rect 45468 17663 45520 17672
rect 45468 17629 45477 17663
rect 45477 17629 45511 17663
rect 45511 17629 45520 17663
rect 45468 17620 45520 17629
rect 45100 17552 45152 17604
rect 45744 17663 45796 17672
rect 45744 17629 45753 17663
rect 45753 17629 45787 17663
rect 45787 17629 45796 17663
rect 46388 17663 46440 17672
rect 45744 17620 45796 17629
rect 46388 17629 46397 17663
rect 46397 17629 46431 17663
rect 46431 17629 46440 17663
rect 46388 17620 46440 17629
rect 46020 17552 46072 17604
rect 46480 17629 46489 17650
rect 46489 17629 46523 17650
rect 46523 17629 46532 17650
rect 46480 17598 46532 17629
rect 47308 17620 47360 17672
rect 47768 17620 47820 17672
rect 49516 17663 49568 17672
rect 38936 17484 38988 17536
rect 39856 17484 39908 17536
rect 40684 17484 40736 17536
rect 42708 17527 42760 17536
rect 42708 17493 42717 17527
rect 42717 17493 42751 17527
rect 42751 17493 42760 17527
rect 42708 17484 42760 17493
rect 46848 17484 46900 17536
rect 47400 17552 47452 17604
rect 48320 17552 48372 17604
rect 49516 17629 49525 17663
rect 49525 17629 49559 17663
rect 49559 17629 49568 17663
rect 49516 17620 49568 17629
rect 49792 17697 49801 17731
rect 49801 17697 49835 17731
rect 49835 17697 49844 17731
rect 52828 17756 52880 17808
rect 52184 17731 52236 17740
rect 49792 17688 49844 17697
rect 50528 17663 50580 17672
rect 50528 17629 50537 17663
rect 50537 17629 50571 17663
rect 50571 17629 50580 17663
rect 50528 17620 50580 17629
rect 52184 17697 52193 17731
rect 52193 17697 52227 17731
rect 52227 17697 52236 17731
rect 52184 17688 52236 17697
rect 52736 17688 52788 17740
rect 50712 17663 50764 17672
rect 50712 17629 50721 17663
rect 50721 17629 50755 17663
rect 50755 17629 50764 17663
rect 50712 17620 50764 17629
rect 51816 17620 51868 17672
rect 52000 17663 52052 17672
rect 52000 17629 52009 17663
rect 52009 17629 52043 17663
rect 52043 17629 52052 17663
rect 52000 17620 52052 17629
rect 52368 17620 52420 17672
rect 53196 17620 53248 17672
rect 55680 17688 55732 17740
rect 55956 17731 56008 17740
rect 55956 17697 55965 17731
rect 55965 17697 55999 17731
rect 55999 17697 56008 17731
rect 55956 17688 56008 17697
rect 56600 17688 56652 17740
rect 53840 17663 53892 17672
rect 53840 17629 53849 17663
rect 53849 17629 53883 17663
rect 53883 17629 53892 17663
rect 53840 17620 53892 17629
rect 54116 17620 54168 17672
rect 55864 17663 55916 17672
rect 55864 17629 55873 17663
rect 55873 17629 55907 17663
rect 55907 17629 55916 17663
rect 55864 17620 55916 17629
rect 50160 17552 50212 17604
rect 50896 17552 50948 17604
rect 47584 17484 47636 17536
rect 48872 17484 48924 17536
rect 51356 17484 51408 17536
rect 51908 17484 51960 17536
rect 54208 17484 54260 17536
rect 54484 17484 54536 17536
rect 54944 17484 54996 17536
rect 57244 17484 57296 17536
rect 57888 17484 57940 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 22100 17280 22152 17332
rect 24768 17280 24820 17332
rect 25504 17280 25556 17332
rect 27712 17280 27764 17332
rect 31208 17323 31260 17332
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 24032 17144 24084 17196
rect 24860 17144 24912 17196
rect 23756 17076 23808 17128
rect 26424 17144 26476 17196
rect 30288 17212 30340 17264
rect 28080 17144 28132 17196
rect 29092 17144 29144 17196
rect 30564 17187 30616 17196
rect 23572 16940 23624 16992
rect 25688 16940 25740 16992
rect 26240 16940 26292 16992
rect 27620 16983 27672 16992
rect 27620 16949 27629 16983
rect 27629 16949 27663 16983
rect 27663 16949 27672 16983
rect 27620 16940 27672 16949
rect 28448 16940 28500 16992
rect 29000 17008 29052 17060
rect 30564 17153 30573 17187
rect 30573 17153 30607 17187
rect 30607 17153 30616 17187
rect 30564 17144 30616 17153
rect 30656 17144 30708 17196
rect 31208 17289 31217 17323
rect 31217 17289 31251 17323
rect 31251 17289 31260 17323
rect 31208 17280 31260 17289
rect 33140 17280 33192 17332
rect 34060 17323 34112 17332
rect 34060 17289 34069 17323
rect 34069 17289 34103 17323
rect 34103 17289 34112 17323
rect 34060 17280 34112 17289
rect 35532 17280 35584 17332
rect 35624 17280 35676 17332
rect 37280 17280 37332 17332
rect 38568 17280 38620 17332
rect 41144 17280 41196 17332
rect 43444 17280 43496 17332
rect 43536 17280 43588 17332
rect 46112 17323 46164 17332
rect 46112 17289 46121 17323
rect 46121 17289 46155 17323
rect 46155 17289 46164 17323
rect 46112 17280 46164 17289
rect 46388 17280 46440 17332
rect 46848 17280 46900 17332
rect 47124 17280 47176 17332
rect 51448 17280 51500 17332
rect 53012 17280 53064 17332
rect 53932 17323 53984 17332
rect 53932 17289 53941 17323
rect 53941 17289 53975 17323
rect 53975 17289 53984 17323
rect 53932 17280 53984 17289
rect 54576 17280 54628 17332
rect 56416 17323 56468 17332
rect 56416 17289 56425 17323
rect 56425 17289 56459 17323
rect 56459 17289 56468 17323
rect 56416 17280 56468 17289
rect 57428 17323 57480 17332
rect 57428 17289 57437 17323
rect 57437 17289 57471 17323
rect 57471 17289 57480 17323
rect 57428 17280 57480 17289
rect 40684 17255 40736 17264
rect 40684 17221 40693 17255
rect 40693 17221 40727 17255
rect 40727 17221 40736 17255
rect 40684 17212 40736 17221
rect 45652 17212 45704 17264
rect 30472 17076 30524 17128
rect 31024 17144 31076 17196
rect 33784 17144 33836 17196
rect 31576 17076 31628 17128
rect 32312 17119 32364 17128
rect 32312 17085 32321 17119
rect 32321 17085 32355 17119
rect 32355 17085 32364 17119
rect 32312 17076 32364 17085
rect 32956 17076 33008 17128
rect 34152 17144 34204 17196
rect 34704 17144 34756 17196
rect 37740 17187 37792 17196
rect 37740 17153 37749 17187
rect 37749 17153 37783 17187
rect 37783 17153 37792 17187
rect 37740 17144 37792 17153
rect 38752 17187 38804 17196
rect 38752 17153 38761 17187
rect 38761 17153 38795 17187
rect 38795 17153 38804 17187
rect 38752 17144 38804 17153
rect 38936 17144 38988 17196
rect 39948 17187 40000 17196
rect 39948 17153 39957 17187
rect 39957 17153 39991 17187
rect 39991 17153 40000 17187
rect 39948 17144 40000 17153
rect 40040 17144 40092 17196
rect 40224 17187 40276 17196
rect 40224 17153 40233 17187
rect 40233 17153 40267 17187
rect 40267 17153 40276 17187
rect 42708 17187 42760 17196
rect 40224 17144 40276 17153
rect 42708 17153 42717 17187
rect 42717 17153 42751 17187
rect 42751 17153 42760 17187
rect 42708 17144 42760 17153
rect 43444 17187 43496 17196
rect 43444 17153 43453 17187
rect 43453 17153 43487 17187
rect 43487 17153 43496 17187
rect 43444 17144 43496 17153
rect 34612 17119 34664 17128
rect 34612 17085 34621 17119
rect 34621 17085 34655 17119
rect 34655 17085 34664 17119
rect 34612 17076 34664 17085
rect 36268 17119 36320 17128
rect 36268 17085 36277 17119
rect 36277 17085 36311 17119
rect 36311 17085 36320 17119
rect 37464 17119 37516 17128
rect 36268 17076 36320 17085
rect 37464 17085 37473 17119
rect 37473 17085 37507 17119
rect 37507 17085 37516 17119
rect 37464 17076 37516 17085
rect 30564 17008 30616 17060
rect 36912 17008 36964 17060
rect 38384 17008 38436 17060
rect 39028 17051 39080 17060
rect 39028 17017 39037 17051
rect 39037 17017 39071 17051
rect 39071 17017 39080 17051
rect 39028 17008 39080 17017
rect 43812 17144 43864 17196
rect 44640 17187 44692 17196
rect 44640 17153 44649 17187
rect 44649 17153 44683 17187
rect 44683 17153 44692 17187
rect 44640 17144 44692 17153
rect 45928 17187 45980 17196
rect 44272 17076 44324 17128
rect 45928 17153 45937 17187
rect 45937 17153 45971 17187
rect 45971 17153 45980 17187
rect 45928 17144 45980 17153
rect 48320 17212 48372 17264
rect 49332 17212 49384 17264
rect 45560 17008 45612 17060
rect 46112 17008 46164 17060
rect 48872 17144 48924 17196
rect 48964 17187 49016 17196
rect 48964 17153 48973 17187
rect 48973 17153 49007 17187
rect 49007 17153 49016 17187
rect 48964 17144 49016 17153
rect 47216 17119 47268 17128
rect 47216 17085 47225 17119
rect 47225 17085 47259 17119
rect 47259 17085 47268 17119
rect 47216 17076 47268 17085
rect 48504 17076 48556 17128
rect 49056 17076 49108 17128
rect 50712 17212 50764 17264
rect 50436 17187 50488 17196
rect 50436 17153 50445 17187
rect 50445 17153 50479 17187
rect 50479 17153 50488 17187
rect 50436 17144 50488 17153
rect 52736 17212 52788 17264
rect 52828 17212 52880 17264
rect 54116 17212 54168 17264
rect 48320 17008 48372 17060
rect 50068 17076 50120 17128
rect 51264 17153 51273 17158
rect 51273 17153 51307 17158
rect 51307 17153 51316 17158
rect 51264 17106 51316 17153
rect 51356 17187 51408 17196
rect 51356 17153 51365 17187
rect 51365 17153 51399 17187
rect 51399 17153 51408 17187
rect 52000 17187 52052 17196
rect 51356 17144 51408 17153
rect 52000 17153 52009 17187
rect 52009 17153 52043 17187
rect 52043 17153 52052 17187
rect 52000 17144 52052 17153
rect 53012 17144 53064 17196
rect 53840 17187 53892 17196
rect 53840 17153 53849 17187
rect 53849 17153 53883 17187
rect 53883 17153 53892 17187
rect 53840 17144 53892 17153
rect 53932 17144 53984 17196
rect 54852 17187 54904 17196
rect 51908 17076 51960 17128
rect 52368 17076 52420 17128
rect 29460 16983 29512 16992
rect 29460 16949 29469 16983
rect 29469 16949 29503 16983
rect 29503 16949 29512 16983
rect 29460 16940 29512 16949
rect 37188 16940 37240 16992
rect 40868 16983 40920 16992
rect 40868 16949 40877 16983
rect 40877 16949 40911 16983
rect 40911 16949 40920 16983
rect 40868 16940 40920 16949
rect 41512 16940 41564 16992
rect 42524 16940 42576 16992
rect 45100 16940 45152 16992
rect 45468 16940 45520 16992
rect 50160 16940 50212 16992
rect 50804 16940 50856 16992
rect 52000 16940 52052 16992
rect 52736 16940 52788 16992
rect 53656 17076 53708 17128
rect 54852 17153 54861 17187
rect 54861 17153 54895 17187
rect 54895 17153 54904 17187
rect 54852 17144 54904 17153
rect 55864 17187 55916 17196
rect 55864 17153 55873 17187
rect 55873 17153 55907 17187
rect 55907 17153 55916 17187
rect 55864 17144 55916 17153
rect 55956 17144 56008 17196
rect 56508 17144 56560 17196
rect 54208 17076 54260 17128
rect 54484 17076 54536 17128
rect 57520 17076 57572 17128
rect 55680 17008 55732 17060
rect 55496 16940 55548 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 23756 16736 23808 16788
rect 29000 16779 29052 16788
rect 29000 16745 29009 16779
rect 29009 16745 29043 16779
rect 29043 16745 29052 16779
rect 29000 16736 29052 16745
rect 30932 16736 30984 16788
rect 31576 16736 31628 16788
rect 26516 16711 26568 16720
rect 26516 16677 26525 16711
rect 26525 16677 26559 16711
rect 26559 16677 26568 16711
rect 26516 16668 26568 16677
rect 27988 16668 28040 16720
rect 29736 16668 29788 16720
rect 22100 16600 22152 16652
rect 23756 16600 23808 16652
rect 26240 16643 26292 16652
rect 26240 16609 26249 16643
rect 26249 16609 26283 16643
rect 26283 16609 26292 16643
rect 26240 16600 26292 16609
rect 27620 16643 27672 16652
rect 27620 16609 27629 16643
rect 27629 16609 27663 16643
rect 27663 16609 27672 16643
rect 27620 16600 27672 16609
rect 30288 16668 30340 16720
rect 32312 16668 32364 16720
rect 36912 16668 36964 16720
rect 33140 16600 33192 16652
rect 38384 16643 38436 16652
rect 26148 16575 26200 16584
rect 26148 16541 26157 16575
rect 26157 16541 26191 16575
rect 26191 16541 26200 16575
rect 26148 16532 26200 16541
rect 26608 16532 26660 16584
rect 23848 16464 23900 16516
rect 24768 16464 24820 16516
rect 25504 16464 25556 16516
rect 28448 16464 28500 16516
rect 29460 16532 29512 16584
rect 30196 16532 30248 16584
rect 30472 16532 30524 16584
rect 31208 16532 31260 16584
rect 29092 16464 29144 16516
rect 33048 16532 33100 16584
rect 33784 16532 33836 16584
rect 34152 16575 34204 16584
rect 34152 16541 34161 16575
rect 34161 16541 34195 16575
rect 34195 16541 34204 16575
rect 34152 16532 34204 16541
rect 36636 16532 36688 16584
rect 26240 16396 26292 16448
rect 26516 16396 26568 16448
rect 27160 16396 27212 16448
rect 32956 16464 33008 16516
rect 34704 16464 34756 16516
rect 30288 16439 30340 16448
rect 30288 16405 30297 16439
rect 30297 16405 30331 16439
rect 30331 16405 30340 16439
rect 30288 16396 30340 16405
rect 31300 16396 31352 16448
rect 32772 16439 32824 16448
rect 32772 16405 32781 16439
rect 32781 16405 32815 16439
rect 32815 16405 32824 16439
rect 32772 16396 32824 16405
rect 33048 16396 33100 16448
rect 34520 16396 34572 16448
rect 38384 16609 38393 16643
rect 38393 16609 38427 16643
rect 38427 16609 38436 16643
rect 38384 16600 38436 16609
rect 37372 16575 37424 16584
rect 37372 16541 37381 16575
rect 37381 16541 37415 16575
rect 37415 16541 37424 16575
rect 37372 16532 37424 16541
rect 38016 16532 38068 16584
rect 38568 16532 38620 16584
rect 38752 16532 38804 16584
rect 39488 16575 39540 16584
rect 39488 16541 39497 16575
rect 39497 16541 39531 16575
rect 39531 16541 39540 16575
rect 40224 16736 40276 16788
rect 42708 16736 42760 16788
rect 45468 16736 45520 16788
rect 47860 16736 47912 16788
rect 39488 16532 39540 16541
rect 40316 16575 40368 16584
rect 40316 16541 40325 16575
rect 40325 16541 40359 16575
rect 40359 16541 40368 16575
rect 40316 16532 40368 16541
rect 41512 16575 41564 16584
rect 41512 16541 41521 16575
rect 41521 16541 41555 16575
rect 41555 16541 41564 16575
rect 41512 16532 41564 16541
rect 41972 16575 42024 16584
rect 41972 16541 41981 16575
rect 41981 16541 42015 16575
rect 42015 16541 42024 16575
rect 41972 16532 42024 16541
rect 44732 16532 44784 16584
rect 46112 16575 46164 16584
rect 46112 16541 46121 16575
rect 46121 16541 46155 16575
rect 46155 16541 46164 16575
rect 46112 16532 46164 16541
rect 46480 16575 46532 16584
rect 37464 16464 37516 16516
rect 42064 16464 42116 16516
rect 43812 16507 43864 16516
rect 43812 16473 43821 16507
rect 43821 16473 43855 16507
rect 43855 16473 43864 16507
rect 43812 16464 43864 16473
rect 45376 16507 45428 16516
rect 45376 16473 45385 16507
rect 45385 16473 45419 16507
rect 45419 16473 45428 16507
rect 45376 16464 45428 16473
rect 37280 16396 37332 16448
rect 37832 16439 37884 16448
rect 37832 16405 37841 16439
rect 37841 16405 37875 16439
rect 37875 16405 37884 16439
rect 37832 16396 37884 16405
rect 38108 16396 38160 16448
rect 40040 16396 40092 16448
rect 46480 16541 46489 16575
rect 46489 16541 46523 16575
rect 46523 16541 46532 16575
rect 46480 16532 46532 16541
rect 46848 16532 46900 16584
rect 47400 16532 47452 16584
rect 46756 16464 46808 16516
rect 48044 16668 48096 16720
rect 48412 16668 48464 16720
rect 50804 16668 50856 16720
rect 52276 16736 52328 16788
rect 53472 16736 53524 16788
rect 53748 16779 53800 16788
rect 53748 16745 53757 16779
rect 53757 16745 53791 16779
rect 53791 16745 53800 16779
rect 53748 16736 53800 16745
rect 54852 16736 54904 16788
rect 56048 16779 56100 16788
rect 56048 16745 56057 16779
rect 56057 16745 56091 16779
rect 56091 16745 56100 16779
rect 56048 16736 56100 16745
rect 56600 16779 56652 16788
rect 56600 16745 56609 16779
rect 56609 16745 56643 16779
rect 56643 16745 56652 16779
rect 56600 16736 56652 16745
rect 47860 16532 47912 16584
rect 48780 16600 48832 16652
rect 53012 16668 53064 16720
rect 50068 16532 50120 16584
rect 50528 16575 50580 16584
rect 50528 16541 50537 16575
rect 50537 16541 50571 16575
rect 50571 16541 50580 16575
rect 50528 16532 50580 16541
rect 50804 16532 50856 16584
rect 51356 16575 51408 16584
rect 51356 16541 51365 16575
rect 51365 16541 51399 16575
rect 51399 16541 51408 16575
rect 51356 16532 51408 16541
rect 52552 16600 52604 16652
rect 53104 16600 53156 16652
rect 52644 16575 52696 16584
rect 48780 16464 48832 16516
rect 49608 16464 49660 16516
rect 48274 16396 48326 16448
rect 48504 16396 48556 16448
rect 50988 16396 51040 16448
rect 51540 16507 51592 16516
rect 51540 16473 51549 16507
rect 51549 16473 51583 16507
rect 51583 16473 51592 16507
rect 51540 16464 51592 16473
rect 52644 16541 52653 16575
rect 52653 16541 52687 16575
rect 52687 16541 52696 16575
rect 52644 16532 52696 16541
rect 53380 16532 53432 16584
rect 53840 16600 53892 16652
rect 56508 16643 56560 16652
rect 54668 16575 54720 16584
rect 54668 16541 54677 16575
rect 54677 16541 54711 16575
rect 54711 16541 54720 16575
rect 54668 16532 54720 16541
rect 55036 16532 55088 16584
rect 55496 16575 55548 16584
rect 55496 16541 55505 16575
rect 55505 16541 55539 16575
rect 55539 16541 55548 16575
rect 55496 16532 55548 16541
rect 55588 16575 55640 16584
rect 55588 16541 55597 16575
rect 55597 16541 55631 16575
rect 55631 16541 55640 16575
rect 55588 16532 55640 16541
rect 56508 16609 56517 16643
rect 56517 16609 56551 16643
rect 56551 16609 56560 16643
rect 56508 16600 56560 16609
rect 52276 16464 52328 16516
rect 53196 16464 53248 16516
rect 54484 16507 54536 16516
rect 54484 16473 54493 16507
rect 54493 16473 54527 16507
rect 54527 16473 54536 16507
rect 54484 16464 54536 16473
rect 56784 16575 56836 16584
rect 56784 16541 56793 16575
rect 56793 16541 56827 16575
rect 56827 16541 56836 16575
rect 56784 16532 56836 16541
rect 52552 16396 52604 16448
rect 53748 16396 53800 16448
rect 56692 16464 56744 16516
rect 56968 16464 57020 16516
rect 56600 16396 56652 16448
rect 57888 16439 57940 16448
rect 57888 16405 57897 16439
rect 57897 16405 57931 16439
rect 57931 16405 57940 16439
rect 57888 16396 57940 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 22100 16192 22152 16244
rect 23572 16192 23624 16244
rect 23756 16235 23808 16244
rect 23756 16201 23765 16235
rect 23765 16201 23799 16235
rect 23799 16201 23808 16235
rect 23756 16192 23808 16201
rect 25504 16235 25556 16244
rect 25504 16201 25513 16235
rect 25513 16201 25547 16235
rect 25547 16201 25556 16235
rect 25504 16192 25556 16201
rect 26148 16192 26200 16244
rect 26608 16235 26660 16244
rect 23848 16124 23900 16176
rect 26608 16201 26617 16235
rect 26617 16201 26651 16235
rect 26651 16201 26660 16235
rect 26608 16192 26660 16201
rect 29000 16192 29052 16244
rect 30564 16192 30616 16244
rect 33048 16192 33100 16244
rect 33692 16192 33744 16244
rect 34428 16192 34480 16244
rect 34704 16235 34756 16244
rect 34704 16201 34713 16235
rect 34713 16201 34747 16235
rect 34747 16201 34756 16235
rect 34704 16192 34756 16201
rect 36820 16235 36872 16244
rect 36820 16201 36829 16235
rect 36829 16201 36863 16235
rect 36863 16201 36872 16235
rect 36820 16192 36872 16201
rect 38108 16235 38160 16244
rect 38108 16201 38117 16235
rect 38117 16201 38151 16235
rect 38151 16201 38160 16235
rect 38108 16192 38160 16201
rect 40224 16192 40276 16244
rect 40868 16192 40920 16244
rect 41144 16235 41196 16244
rect 41144 16201 41153 16235
rect 41153 16201 41187 16235
rect 41187 16201 41196 16235
rect 41144 16192 41196 16201
rect 41420 16192 41472 16244
rect 42800 16235 42852 16244
rect 42800 16201 42809 16235
rect 42809 16201 42843 16235
rect 42843 16201 42852 16235
rect 42800 16192 42852 16201
rect 43812 16192 43864 16244
rect 44732 16235 44784 16244
rect 44732 16201 44741 16235
rect 44741 16201 44775 16235
rect 44775 16201 44784 16235
rect 44732 16192 44784 16201
rect 46204 16235 46256 16244
rect 46204 16201 46213 16235
rect 46213 16201 46247 16235
rect 46247 16201 46256 16235
rect 46204 16192 46256 16201
rect 30472 16124 30524 16176
rect 31208 16124 31260 16176
rect 26056 16056 26108 16108
rect 26424 16099 26476 16108
rect 26424 16065 26433 16099
rect 26433 16065 26467 16099
rect 26467 16065 26476 16099
rect 26424 16056 26476 16065
rect 27436 16099 27488 16108
rect 27436 16065 27445 16099
rect 27445 16065 27479 16099
rect 27479 16065 27488 16099
rect 27436 16056 27488 16065
rect 29736 16099 29788 16108
rect 29736 16065 29745 16099
rect 29745 16065 29779 16099
rect 29779 16065 29788 16099
rect 29736 16056 29788 16065
rect 29920 16099 29972 16108
rect 29920 16065 29929 16099
rect 29929 16065 29963 16099
rect 29963 16065 29972 16099
rect 29920 16056 29972 16065
rect 30196 16056 30248 16108
rect 31024 16099 31076 16108
rect 31024 16065 31033 16099
rect 31033 16065 31067 16099
rect 31067 16065 31076 16099
rect 31024 16056 31076 16065
rect 31300 16099 31352 16108
rect 25044 15988 25096 16040
rect 26148 16031 26200 16040
rect 26148 15997 26157 16031
rect 26157 15997 26191 16031
rect 26191 15997 26200 16031
rect 26148 15988 26200 15997
rect 26332 16031 26384 16040
rect 26332 15997 26341 16031
rect 26341 15997 26375 16031
rect 26375 15997 26384 16031
rect 27160 16031 27212 16040
rect 26332 15988 26384 15997
rect 27160 15997 27169 16031
rect 27169 15997 27203 16031
rect 27203 15997 27212 16031
rect 27160 15988 27212 15997
rect 31300 16065 31309 16099
rect 31309 16065 31343 16099
rect 31343 16065 31352 16099
rect 31300 16056 31352 16065
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 33416 16056 33468 16108
rect 32772 16031 32824 16040
rect 32772 15997 32781 16031
rect 32781 15997 32815 16031
rect 32815 15997 32824 16031
rect 32772 15988 32824 15997
rect 33324 15988 33376 16040
rect 35440 15988 35492 16040
rect 35624 16031 35676 16040
rect 35624 15997 35633 16031
rect 35633 15997 35667 16031
rect 35667 15997 35676 16031
rect 35624 15988 35676 15997
rect 26976 15920 27028 15972
rect 27896 15920 27948 15972
rect 31116 15920 31168 15972
rect 32496 15920 32548 15972
rect 36728 16099 36780 16108
rect 36728 16065 36737 16099
rect 36737 16065 36771 16099
rect 36771 16065 36780 16099
rect 36728 16056 36780 16065
rect 37648 16056 37700 16108
rect 38016 16099 38068 16108
rect 38016 16065 38025 16099
rect 38025 16065 38059 16099
rect 38059 16065 38068 16099
rect 38016 16056 38068 16065
rect 38752 16056 38804 16108
rect 40040 16056 40092 16108
rect 41512 16099 41564 16108
rect 39948 15988 40000 16040
rect 41512 16065 41521 16099
rect 41521 16065 41555 16099
rect 41555 16065 41564 16099
rect 41512 16056 41564 16065
rect 41972 16056 42024 16108
rect 42708 16099 42760 16108
rect 42708 16065 42717 16099
rect 42717 16065 42751 16099
rect 42751 16065 42760 16099
rect 42708 16056 42760 16065
rect 45192 16124 45244 16176
rect 47216 16192 47268 16244
rect 48504 16235 48556 16244
rect 47860 16124 47912 16176
rect 48504 16201 48513 16235
rect 48513 16201 48547 16235
rect 48547 16201 48556 16235
rect 48504 16192 48556 16201
rect 49240 16192 49292 16244
rect 49976 16192 50028 16244
rect 50804 16192 50856 16244
rect 50988 16192 51040 16244
rect 51540 16192 51592 16244
rect 54116 16192 54168 16244
rect 54484 16192 54536 16244
rect 55680 16192 55732 16244
rect 56508 16192 56560 16244
rect 45560 16099 45612 16108
rect 42524 15988 42576 16040
rect 44088 15988 44140 16040
rect 44456 15988 44508 16040
rect 45560 16065 45569 16099
rect 45569 16065 45603 16099
rect 45603 16065 45612 16099
rect 45560 16056 45612 16065
rect 45744 16099 45796 16108
rect 45744 16065 45752 16099
rect 45752 16065 45786 16099
rect 45786 16065 45796 16099
rect 45744 16056 45796 16065
rect 46020 16056 46072 16108
rect 45836 16031 45888 16040
rect 45836 15997 45845 16031
rect 45845 15997 45879 16031
rect 45879 15997 45888 16031
rect 45836 15988 45888 15997
rect 46204 16056 46256 16108
rect 46848 16056 46900 16108
rect 46664 15988 46716 16040
rect 47400 16056 47452 16108
rect 48136 16056 48188 16108
rect 48688 16099 48740 16108
rect 48688 16065 48697 16099
rect 48697 16065 48731 16099
rect 48731 16065 48740 16099
rect 48688 16056 48740 16065
rect 50160 16056 50212 16108
rect 43628 15963 43680 15972
rect 43628 15929 43637 15963
rect 43637 15929 43671 15963
rect 43671 15929 43680 15963
rect 43628 15920 43680 15929
rect 26332 15852 26384 15904
rect 28448 15852 28500 15904
rect 29460 15852 29512 15904
rect 37832 15852 37884 15904
rect 41604 15852 41656 15904
rect 46756 15920 46808 15972
rect 46112 15852 46164 15904
rect 47032 15988 47084 16040
rect 47952 15963 48004 15972
rect 47952 15929 47961 15963
rect 47961 15929 47995 15963
rect 47995 15929 48004 15963
rect 47952 15920 48004 15929
rect 48964 16031 49016 16040
rect 48964 15997 48973 16031
rect 48973 15997 49007 16031
rect 49007 15997 49016 16031
rect 48964 15988 49016 15997
rect 49976 15988 50028 16040
rect 50436 16056 50488 16108
rect 50620 16099 50672 16108
rect 50620 16065 50629 16099
rect 50629 16065 50663 16099
rect 50663 16065 50672 16099
rect 50620 16056 50672 16065
rect 50804 16099 50856 16108
rect 50804 16065 50813 16099
rect 50813 16065 50847 16099
rect 50847 16065 50856 16099
rect 50804 16056 50856 16065
rect 51172 16124 51224 16176
rect 51356 16031 51408 16040
rect 51356 15997 51365 16031
rect 51365 15997 51399 16031
rect 51399 15997 51408 16031
rect 51356 15988 51408 15997
rect 51540 16099 51592 16108
rect 51540 16065 51549 16099
rect 51549 16065 51583 16099
rect 51583 16065 51592 16099
rect 51540 16056 51592 16065
rect 52000 16056 52052 16108
rect 53840 16099 53892 16108
rect 53840 16065 53849 16099
rect 53849 16065 53883 16099
rect 53883 16065 53892 16099
rect 53840 16056 53892 16065
rect 53748 15988 53800 16040
rect 49424 15920 49476 15972
rect 49700 15920 49752 15972
rect 48964 15852 49016 15904
rect 50252 15852 50304 15904
rect 51080 15920 51132 15972
rect 54208 15988 54260 16040
rect 55220 16056 55272 16108
rect 55588 16056 55640 16108
rect 55496 15988 55548 16040
rect 54484 15920 54536 15972
rect 54852 15920 54904 15972
rect 51448 15852 51500 15904
rect 55128 15852 55180 15904
rect 56600 15895 56652 15904
rect 56600 15861 56609 15895
rect 56609 15861 56643 15895
rect 56643 15861 56652 15895
rect 56600 15852 56652 15861
rect 57152 15895 57204 15904
rect 57152 15861 57161 15895
rect 57161 15861 57195 15895
rect 57195 15861 57204 15895
rect 57152 15852 57204 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 23572 15648 23624 15700
rect 24952 15648 25004 15700
rect 25412 15691 25464 15700
rect 25412 15657 25421 15691
rect 25421 15657 25455 15691
rect 25455 15657 25464 15691
rect 25412 15648 25464 15657
rect 26056 15648 26108 15700
rect 27436 15648 27488 15700
rect 28080 15648 28132 15700
rect 30840 15648 30892 15700
rect 31208 15648 31260 15700
rect 32772 15648 32824 15700
rect 35624 15691 35676 15700
rect 35624 15657 35633 15691
rect 35633 15657 35667 15691
rect 35667 15657 35676 15691
rect 35624 15648 35676 15657
rect 36268 15648 36320 15700
rect 37648 15691 37700 15700
rect 37648 15657 37657 15691
rect 37657 15657 37691 15691
rect 37691 15657 37700 15691
rect 37648 15648 37700 15657
rect 38476 15691 38528 15700
rect 38476 15657 38485 15691
rect 38485 15657 38519 15691
rect 38519 15657 38528 15691
rect 38476 15648 38528 15657
rect 45744 15648 45796 15700
rect 45836 15648 45888 15700
rect 24032 15580 24084 15632
rect 26516 15580 26568 15632
rect 27896 15623 27948 15632
rect 27896 15589 27905 15623
rect 27905 15589 27939 15623
rect 27939 15589 27948 15623
rect 27896 15580 27948 15589
rect 28816 15580 28868 15632
rect 22560 15512 22612 15564
rect 24308 15512 24360 15564
rect 29920 15580 29972 15632
rect 36728 15580 36780 15632
rect 42800 15580 42852 15632
rect 44180 15580 44232 15632
rect 44364 15580 44416 15632
rect 44824 15580 44876 15632
rect 47400 15648 47452 15700
rect 29828 15555 29880 15564
rect 29828 15521 29837 15555
rect 29837 15521 29871 15555
rect 29871 15521 29880 15555
rect 29828 15512 29880 15521
rect 22836 15444 22888 15496
rect 23572 15487 23624 15496
rect 23572 15453 23581 15487
rect 23581 15453 23615 15487
rect 23615 15453 23624 15487
rect 23572 15444 23624 15453
rect 23756 15444 23808 15496
rect 26240 15444 26292 15496
rect 27988 15444 28040 15496
rect 28540 15444 28592 15496
rect 28724 15487 28776 15496
rect 28724 15453 28733 15487
rect 28733 15453 28767 15487
rect 28767 15453 28776 15487
rect 28724 15444 28776 15453
rect 29000 15487 29052 15496
rect 27068 15376 27120 15428
rect 27528 15419 27580 15428
rect 27528 15385 27537 15419
rect 27537 15385 27571 15419
rect 27571 15385 27580 15419
rect 27528 15376 27580 15385
rect 29000 15453 29009 15487
rect 29009 15453 29043 15487
rect 29043 15453 29052 15487
rect 29000 15444 29052 15453
rect 30196 15444 30248 15496
rect 30840 15444 30892 15496
rect 31392 15444 31444 15496
rect 32220 15444 32272 15496
rect 32956 15487 33008 15496
rect 32956 15453 32965 15487
rect 32965 15453 32999 15487
rect 32999 15453 33008 15487
rect 32956 15444 33008 15453
rect 33324 15444 33376 15496
rect 34152 15444 34204 15496
rect 30932 15376 30984 15428
rect 31024 15419 31076 15428
rect 31024 15385 31033 15419
rect 31033 15385 31067 15419
rect 31067 15385 31076 15419
rect 32312 15419 32364 15428
rect 31024 15376 31076 15385
rect 32312 15385 32321 15419
rect 32321 15385 32355 15419
rect 32355 15385 32364 15419
rect 32312 15376 32364 15385
rect 34796 15376 34848 15428
rect 22376 15308 22428 15360
rect 23296 15308 23348 15360
rect 28632 15308 28684 15360
rect 28908 15308 28960 15360
rect 31300 15308 31352 15360
rect 33416 15308 33468 15360
rect 34336 15351 34388 15360
rect 34336 15317 34345 15351
rect 34345 15317 34379 15351
rect 34379 15317 34388 15351
rect 34336 15308 34388 15317
rect 34704 15308 34756 15360
rect 35900 15444 35952 15496
rect 36360 15512 36412 15564
rect 39028 15555 39080 15564
rect 39028 15521 39037 15555
rect 39037 15521 39071 15555
rect 39071 15521 39080 15555
rect 39028 15512 39080 15521
rect 45376 15555 45428 15564
rect 45376 15521 45385 15555
rect 45385 15521 45419 15555
rect 45419 15521 45428 15555
rect 45376 15512 45428 15521
rect 36636 15487 36688 15496
rect 36636 15453 36645 15487
rect 36645 15453 36679 15487
rect 36679 15453 36688 15487
rect 36636 15444 36688 15453
rect 36360 15419 36412 15428
rect 36360 15385 36369 15419
rect 36369 15385 36403 15419
rect 36403 15385 36412 15419
rect 36360 15376 36412 15385
rect 36452 15419 36504 15428
rect 36452 15385 36461 15419
rect 36461 15385 36495 15419
rect 36495 15385 36504 15419
rect 36452 15376 36504 15385
rect 37832 15444 37884 15496
rect 39120 15444 39172 15496
rect 38660 15376 38712 15428
rect 39948 15376 40000 15428
rect 42524 15376 42576 15428
rect 43260 15444 43312 15496
rect 43628 15376 43680 15428
rect 46112 15512 46164 15564
rect 47952 15580 48004 15632
rect 46664 15512 46716 15564
rect 47400 15555 47452 15564
rect 47400 15521 47409 15555
rect 47409 15521 47443 15555
rect 47443 15521 47452 15555
rect 47400 15512 47452 15521
rect 47492 15555 47544 15564
rect 47492 15521 47501 15555
rect 47501 15521 47535 15555
rect 47535 15521 47544 15555
rect 47492 15512 47544 15521
rect 47768 15512 47820 15564
rect 48688 15648 48740 15700
rect 50160 15648 50212 15700
rect 50620 15648 50672 15700
rect 51632 15648 51684 15700
rect 54944 15691 54996 15700
rect 54944 15657 54953 15691
rect 54953 15657 54987 15691
rect 54987 15657 54996 15691
rect 54944 15648 54996 15657
rect 57520 15691 57572 15700
rect 57520 15657 57529 15691
rect 57529 15657 57563 15691
rect 57563 15657 57572 15691
rect 57520 15648 57572 15657
rect 50068 15580 50120 15632
rect 51816 15580 51868 15632
rect 51908 15512 51960 15564
rect 56784 15580 56836 15632
rect 46848 15444 46900 15496
rect 47032 15444 47084 15496
rect 47584 15487 47636 15496
rect 47584 15453 47593 15487
rect 47593 15453 47627 15487
rect 47627 15453 47636 15487
rect 47584 15444 47636 15453
rect 48228 15444 48280 15496
rect 50712 15444 50764 15496
rect 52276 15487 52328 15496
rect 47400 15376 47452 15428
rect 38752 15308 38804 15360
rect 39396 15308 39448 15360
rect 40868 15308 40920 15360
rect 45284 15351 45336 15360
rect 45284 15317 45293 15351
rect 45293 15317 45327 15351
rect 45327 15317 45336 15351
rect 45284 15308 45336 15317
rect 45652 15308 45704 15360
rect 45744 15308 45796 15360
rect 46204 15308 46256 15360
rect 46756 15308 46808 15360
rect 47860 15351 47912 15360
rect 47860 15317 47869 15351
rect 47869 15317 47903 15351
rect 47903 15317 47912 15351
rect 47860 15308 47912 15317
rect 49240 15376 49292 15428
rect 49976 15376 50028 15428
rect 52276 15453 52285 15487
rect 52285 15453 52319 15487
rect 52319 15453 52328 15487
rect 52276 15444 52328 15453
rect 52460 15444 52512 15496
rect 53196 15487 53248 15496
rect 53196 15453 53205 15487
rect 53205 15453 53239 15487
rect 53239 15453 53248 15487
rect 53196 15444 53248 15453
rect 53472 15444 53524 15496
rect 52920 15376 52972 15428
rect 56600 15512 56652 15564
rect 55220 15444 55272 15496
rect 56692 15444 56744 15496
rect 54484 15376 54536 15428
rect 57152 15376 57204 15428
rect 49516 15308 49568 15360
rect 52828 15351 52880 15360
rect 52828 15317 52837 15351
rect 52837 15317 52871 15351
rect 52871 15317 52880 15351
rect 52828 15308 52880 15317
rect 53656 15308 53708 15360
rect 53840 15308 53892 15360
rect 56232 15308 56284 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 23572 15104 23624 15156
rect 24032 15147 24084 15156
rect 24032 15113 24041 15147
rect 24041 15113 24075 15147
rect 24075 15113 24084 15147
rect 24032 15104 24084 15113
rect 24768 15104 24820 15156
rect 26424 15104 26476 15156
rect 29000 15104 29052 15156
rect 29644 15104 29696 15156
rect 22836 15079 22888 15088
rect 22836 15045 22845 15079
rect 22845 15045 22879 15079
rect 22879 15045 22888 15079
rect 26516 15079 26568 15088
rect 22836 15036 22888 15045
rect 26516 15045 26525 15079
rect 26525 15045 26559 15079
rect 26559 15045 26568 15079
rect 26516 15036 26568 15045
rect 26976 15036 27028 15088
rect 29920 15036 29972 15088
rect 31116 15036 31168 15088
rect 31392 15036 31444 15088
rect 34428 15036 34480 15088
rect 21364 14968 21416 15020
rect 25504 14968 25556 15020
rect 24124 14943 24176 14952
rect 24124 14909 24133 14943
rect 24133 14909 24167 14943
rect 24167 14909 24176 14943
rect 24124 14900 24176 14909
rect 24308 14943 24360 14952
rect 24308 14909 24317 14943
rect 24317 14909 24351 14943
rect 24351 14909 24360 14943
rect 24308 14900 24360 14909
rect 24768 14900 24820 14952
rect 27068 14968 27120 15020
rect 27620 15011 27672 15020
rect 27620 14977 27629 15011
rect 27629 14977 27663 15011
rect 27663 14977 27672 15011
rect 27620 14968 27672 14977
rect 27988 14968 28040 15020
rect 28816 14968 28868 15020
rect 30012 15011 30064 15020
rect 30012 14977 30021 15011
rect 30021 14977 30055 15011
rect 30055 14977 30064 15011
rect 30012 14968 30064 14977
rect 30104 14968 30156 15020
rect 30932 14968 30984 15020
rect 29184 14943 29236 14952
rect 29184 14909 29193 14943
rect 29193 14909 29227 14943
rect 29227 14909 29236 14943
rect 29184 14900 29236 14909
rect 31852 14968 31904 15020
rect 32220 14968 32272 15020
rect 34336 14968 34388 15020
rect 36176 15104 36228 15156
rect 36636 15104 36688 15156
rect 37372 15104 37424 15156
rect 39028 15104 39080 15156
rect 41972 15104 42024 15156
rect 43444 15104 43496 15156
rect 43720 15104 43772 15156
rect 44180 15104 44232 15156
rect 44640 15147 44692 15156
rect 44640 15113 44649 15147
rect 44649 15113 44683 15147
rect 44683 15113 44692 15147
rect 44640 15104 44692 15113
rect 45192 15104 45244 15156
rect 45928 15104 45980 15156
rect 47860 15104 47912 15156
rect 48504 15104 48556 15156
rect 35348 15011 35400 15020
rect 35348 14977 35357 15011
rect 35357 14977 35391 15011
rect 35391 14977 35400 15011
rect 35348 14968 35400 14977
rect 39120 15036 39172 15088
rect 36360 15011 36412 15020
rect 36360 14977 36369 15011
rect 36369 14977 36403 15011
rect 36403 14977 36412 15011
rect 36360 14968 36412 14977
rect 36544 15011 36596 15020
rect 36544 14977 36553 15011
rect 36553 14977 36587 15011
rect 36587 14977 36596 15011
rect 36544 14968 36596 14977
rect 37924 14968 37976 15020
rect 39304 15011 39356 15020
rect 39304 14977 39313 15011
rect 39313 14977 39347 15011
rect 39347 14977 39356 15011
rect 39948 15036 40000 15088
rect 41420 15036 41472 15088
rect 39304 14968 39356 14977
rect 43536 15011 43588 15020
rect 43536 14977 43545 15011
rect 43545 14977 43579 15011
rect 43579 14977 43588 15011
rect 43536 14968 43588 14977
rect 28908 14832 28960 14884
rect 21364 14807 21416 14816
rect 21364 14773 21373 14807
rect 21373 14773 21407 14807
rect 21407 14773 21416 14807
rect 21364 14764 21416 14773
rect 27528 14764 27580 14816
rect 28264 14807 28316 14816
rect 28264 14773 28273 14807
rect 28273 14773 28307 14807
rect 28307 14773 28316 14807
rect 28264 14764 28316 14773
rect 30196 14764 30248 14816
rect 32312 14900 32364 14952
rect 32680 14900 32732 14952
rect 35624 14900 35676 14952
rect 32496 14832 32548 14884
rect 32588 14832 32640 14884
rect 35808 14832 35860 14884
rect 37740 14900 37792 14952
rect 38292 14900 38344 14952
rect 39120 14943 39172 14952
rect 39120 14909 39129 14943
rect 39129 14909 39163 14943
rect 39163 14909 39172 14943
rect 39120 14900 39172 14909
rect 31760 14764 31812 14816
rect 32864 14764 32916 14816
rect 34704 14764 34756 14816
rect 37464 14807 37516 14816
rect 37464 14773 37473 14807
rect 37473 14773 37507 14807
rect 37507 14773 37516 14807
rect 37464 14764 37516 14773
rect 38200 14764 38252 14816
rect 38844 14832 38896 14884
rect 39488 14900 39540 14952
rect 43720 15011 43772 15020
rect 43720 14977 43729 15011
rect 43729 14977 43763 15011
rect 43763 14977 43772 15011
rect 44824 15011 44876 15020
rect 43720 14968 43772 14977
rect 44824 14977 44833 15011
rect 44833 14977 44867 15011
rect 44867 14977 44876 15011
rect 44824 14968 44876 14977
rect 44916 15011 44968 15020
rect 44916 14977 44925 15011
rect 44925 14977 44959 15011
rect 44959 14977 44968 15011
rect 44916 14968 44968 14977
rect 45192 14968 45244 15020
rect 45652 15011 45704 15020
rect 45652 14977 45661 15011
rect 45661 14977 45695 15011
rect 45695 14977 45704 15011
rect 45652 14968 45704 14977
rect 45744 15011 45796 15020
rect 45744 14977 45753 15011
rect 45753 14977 45787 15011
rect 45787 14977 45796 15011
rect 45928 15011 45980 15020
rect 45744 14968 45796 14977
rect 45928 14977 45937 15011
rect 45937 14977 45971 15011
rect 45971 14977 45980 15011
rect 45928 14968 45980 14977
rect 46204 15036 46256 15088
rect 46112 14968 46164 15020
rect 47400 15036 47452 15088
rect 47768 15079 47820 15088
rect 47768 15045 47777 15079
rect 47777 15045 47811 15079
rect 47811 15045 47820 15079
rect 47768 15036 47820 15045
rect 49792 15104 49844 15156
rect 48044 14968 48096 15020
rect 48780 15011 48832 15020
rect 48780 14977 48789 15011
rect 48789 14977 48823 15011
rect 48823 14977 48832 15011
rect 48780 14968 48832 14977
rect 43904 14875 43956 14884
rect 43904 14841 43913 14875
rect 43913 14841 43947 14875
rect 43947 14841 43956 14875
rect 43904 14832 43956 14841
rect 39212 14764 39264 14816
rect 43812 14764 43864 14816
rect 44548 14900 44600 14952
rect 46664 14900 46716 14952
rect 48688 14900 48740 14952
rect 48872 14943 48924 14952
rect 48872 14909 48881 14943
rect 48881 14909 48915 14943
rect 48915 14909 48924 14943
rect 48872 14900 48924 14909
rect 45468 14832 45520 14884
rect 45560 14832 45612 14884
rect 48412 14832 48464 14884
rect 48504 14832 48556 14884
rect 49332 14968 49384 15020
rect 49332 14832 49384 14884
rect 49976 15104 50028 15156
rect 51448 15104 51500 15156
rect 51264 15036 51316 15088
rect 50252 14968 50304 15020
rect 50344 15011 50396 15020
rect 50344 14977 50353 15011
rect 50353 14977 50387 15011
rect 50387 14977 50396 15011
rect 50896 15011 50948 15020
rect 50344 14968 50396 14977
rect 50068 14943 50120 14952
rect 50068 14909 50077 14943
rect 50077 14909 50111 14943
rect 50111 14909 50120 14943
rect 50896 14977 50905 15011
rect 50905 14977 50939 15011
rect 50939 14977 50948 15011
rect 50896 14968 50948 14977
rect 51448 14968 51500 15020
rect 51724 14968 51776 15020
rect 53288 15147 53340 15156
rect 53288 15113 53297 15147
rect 53297 15113 53331 15147
rect 53331 15113 53340 15147
rect 53288 15104 53340 15113
rect 54576 15104 54628 15156
rect 52828 15036 52880 15088
rect 53012 15036 53064 15088
rect 54668 15036 54720 15088
rect 54024 15011 54076 15020
rect 50068 14900 50120 14909
rect 51632 14900 51684 14952
rect 45928 14764 45980 14816
rect 47032 14764 47084 14816
rect 47216 14764 47268 14816
rect 48228 14764 48280 14816
rect 50620 14764 50672 14816
rect 51080 14764 51132 14816
rect 54024 14977 54033 15011
rect 54033 14977 54067 15011
rect 54067 14977 54076 15011
rect 54024 14968 54076 14977
rect 53288 14900 53340 14952
rect 54208 14968 54260 15020
rect 54392 15011 54444 15020
rect 54392 14977 54401 15011
rect 54401 14977 54435 15011
rect 54435 14977 54444 15011
rect 55220 15011 55272 15020
rect 54392 14968 54444 14977
rect 55220 14977 55229 15011
rect 55229 14977 55263 15011
rect 55263 14977 55272 15011
rect 55220 14968 55272 14977
rect 55496 15011 55548 15020
rect 55496 14977 55505 15011
rect 55505 14977 55539 15011
rect 55539 14977 55548 15011
rect 55496 14968 55548 14977
rect 55588 14968 55640 15020
rect 55956 14968 56008 15020
rect 56968 15011 57020 15020
rect 56968 14977 56977 15011
rect 56977 14977 57011 15011
rect 57011 14977 57020 15011
rect 56968 14968 57020 14977
rect 52276 14832 52328 14884
rect 53472 14832 53524 14884
rect 54116 14832 54168 14884
rect 55680 14832 55732 14884
rect 57888 14764 57940 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 24124 14560 24176 14612
rect 26240 14560 26292 14612
rect 27620 14560 27672 14612
rect 28540 14560 28592 14612
rect 29920 14560 29972 14612
rect 32312 14560 32364 14612
rect 32404 14560 32456 14612
rect 33416 14603 33468 14612
rect 33416 14569 33425 14603
rect 33425 14569 33459 14603
rect 33459 14569 33468 14603
rect 33416 14560 33468 14569
rect 35440 14560 35492 14612
rect 36544 14603 36596 14612
rect 36544 14569 36553 14603
rect 36553 14569 36587 14603
rect 36587 14569 36596 14603
rect 36544 14560 36596 14569
rect 37924 14603 37976 14612
rect 22376 14399 22428 14408
rect 22376 14365 22385 14399
rect 22385 14365 22419 14399
rect 22419 14365 22428 14399
rect 22376 14356 22428 14365
rect 23296 14399 23348 14408
rect 23296 14365 23305 14399
rect 23305 14365 23339 14399
rect 23339 14365 23348 14399
rect 23296 14356 23348 14365
rect 24676 14356 24728 14408
rect 24952 14331 25004 14340
rect 24952 14297 24961 14331
rect 24961 14297 24995 14331
rect 24995 14297 25004 14331
rect 24952 14288 25004 14297
rect 29092 14492 29144 14544
rect 32680 14492 32732 14544
rect 27712 14424 27764 14476
rect 28172 14424 28224 14476
rect 28264 14424 28316 14476
rect 26516 14331 26568 14340
rect 26516 14297 26525 14331
rect 26525 14297 26559 14331
rect 26559 14297 26568 14331
rect 27620 14356 27672 14408
rect 31116 14356 31168 14408
rect 31392 14399 31444 14408
rect 31392 14365 31401 14399
rect 31401 14365 31435 14399
rect 31435 14365 31444 14399
rect 31392 14356 31444 14365
rect 31576 14399 31628 14408
rect 31576 14365 31585 14399
rect 31585 14365 31619 14399
rect 31619 14365 31628 14399
rect 32312 14399 32364 14408
rect 31576 14356 31628 14365
rect 32312 14365 32321 14399
rect 32321 14365 32355 14399
rect 32355 14365 32364 14399
rect 32312 14356 32364 14365
rect 32496 14399 32548 14408
rect 32496 14365 32505 14399
rect 32505 14365 32539 14399
rect 32539 14365 32548 14399
rect 32496 14356 32548 14365
rect 32588 14399 32640 14408
rect 32588 14365 32597 14399
rect 32597 14365 32631 14399
rect 32631 14365 32640 14399
rect 32588 14356 32640 14365
rect 32864 14356 32916 14408
rect 26516 14288 26568 14297
rect 26148 14220 26200 14272
rect 28264 14288 28316 14340
rect 27896 14220 27948 14272
rect 29552 14288 29604 14340
rect 33784 14424 33836 14476
rect 36268 14492 36320 14544
rect 37924 14569 37933 14603
rect 37933 14569 37967 14603
rect 37967 14569 37976 14603
rect 37924 14560 37976 14569
rect 38384 14603 38436 14612
rect 38384 14569 38393 14603
rect 38393 14569 38427 14603
rect 38427 14569 38436 14603
rect 38384 14560 38436 14569
rect 40592 14603 40644 14612
rect 40592 14569 40601 14603
rect 40601 14569 40635 14603
rect 40635 14569 40644 14603
rect 40592 14560 40644 14569
rect 41420 14603 41472 14612
rect 41420 14569 41429 14603
rect 41429 14569 41463 14603
rect 41463 14569 41472 14603
rect 41420 14560 41472 14569
rect 36820 14492 36872 14544
rect 39488 14492 39540 14544
rect 34888 14399 34940 14408
rect 33600 14288 33652 14340
rect 34888 14365 34897 14399
rect 34897 14365 34931 14399
rect 34931 14365 34940 14399
rect 34888 14356 34940 14365
rect 35348 14424 35400 14476
rect 36360 14424 36412 14476
rect 39304 14424 39356 14476
rect 40592 14424 40644 14476
rect 37556 14399 37608 14408
rect 37556 14365 37565 14399
rect 37565 14365 37599 14399
rect 37599 14365 37608 14399
rect 37556 14356 37608 14365
rect 28908 14263 28960 14272
rect 28908 14229 28917 14263
rect 28917 14229 28951 14263
rect 28951 14229 28960 14263
rect 28908 14220 28960 14229
rect 33876 14220 33928 14272
rect 33968 14220 34020 14272
rect 34428 14220 34480 14272
rect 37004 14288 37056 14340
rect 38384 14356 38436 14408
rect 38660 14356 38712 14408
rect 38476 14288 38528 14340
rect 39948 14356 40000 14408
rect 41696 14356 41748 14408
rect 43076 14560 43128 14612
rect 43260 14492 43312 14544
rect 44916 14560 44968 14612
rect 44180 14492 44232 14544
rect 45560 14560 45612 14612
rect 45652 14603 45704 14612
rect 45652 14569 45661 14603
rect 45661 14569 45695 14603
rect 45695 14569 45704 14603
rect 45652 14560 45704 14569
rect 46020 14560 46072 14612
rect 46940 14560 46992 14612
rect 48044 14603 48096 14612
rect 48044 14569 48053 14603
rect 48053 14569 48087 14603
rect 48087 14569 48096 14603
rect 48044 14560 48096 14569
rect 45836 14492 45888 14544
rect 42524 14399 42576 14408
rect 42524 14365 42533 14399
rect 42533 14365 42567 14399
rect 42567 14365 42576 14399
rect 42524 14356 42576 14365
rect 43904 14356 43956 14408
rect 45652 14356 45704 14408
rect 46296 14492 46348 14544
rect 48688 14492 48740 14544
rect 48872 14560 48924 14612
rect 50620 14560 50672 14612
rect 51172 14603 51224 14612
rect 51172 14569 51181 14603
rect 51181 14569 51215 14603
rect 51215 14569 51224 14603
rect 51172 14560 51224 14569
rect 51908 14560 51960 14612
rect 52184 14560 52236 14612
rect 52552 14603 52604 14612
rect 52552 14569 52561 14603
rect 52561 14569 52595 14603
rect 52595 14569 52604 14603
rect 52552 14560 52604 14569
rect 52920 14560 52972 14612
rect 54392 14603 54444 14612
rect 54392 14569 54401 14603
rect 54401 14569 54435 14603
rect 54435 14569 54444 14603
rect 54392 14560 54444 14569
rect 55128 14560 55180 14612
rect 56232 14603 56284 14612
rect 56232 14569 56241 14603
rect 56241 14569 56275 14603
rect 56275 14569 56284 14603
rect 56232 14560 56284 14569
rect 57612 14560 57664 14612
rect 49792 14535 49844 14544
rect 49792 14501 49801 14535
rect 49801 14501 49835 14535
rect 49835 14501 49844 14535
rect 49792 14492 49844 14501
rect 46664 14424 46716 14476
rect 47032 14399 47084 14408
rect 44180 14288 44232 14340
rect 45376 14288 45428 14340
rect 36176 14220 36228 14272
rect 36728 14263 36780 14272
rect 36728 14229 36755 14263
rect 36755 14229 36780 14263
rect 36728 14220 36780 14229
rect 38200 14220 38252 14272
rect 41972 14220 42024 14272
rect 43444 14220 43496 14272
rect 45560 14220 45612 14272
rect 45744 14220 45796 14272
rect 47032 14365 47041 14399
rect 47041 14365 47075 14399
rect 47075 14365 47084 14399
rect 47032 14356 47084 14365
rect 47124 14399 47176 14408
rect 47124 14365 47133 14399
rect 47133 14365 47167 14399
rect 47167 14365 47176 14399
rect 47400 14399 47452 14408
rect 47124 14356 47176 14365
rect 47400 14365 47409 14399
rect 47409 14365 47443 14399
rect 47443 14365 47452 14399
rect 47400 14356 47452 14365
rect 46940 14288 46992 14340
rect 47768 14288 47820 14340
rect 48412 14356 48464 14408
rect 48688 14356 48740 14408
rect 49056 14356 49108 14408
rect 49976 14424 50028 14476
rect 49332 14356 49384 14408
rect 50160 14492 50212 14544
rect 53104 14492 53156 14544
rect 52644 14424 52696 14476
rect 51172 14356 51224 14408
rect 51908 14399 51960 14408
rect 51908 14365 51917 14399
rect 51917 14365 51951 14399
rect 51951 14365 51960 14399
rect 51908 14356 51960 14365
rect 52092 14399 52144 14408
rect 52092 14365 52101 14399
rect 52101 14365 52135 14399
rect 52135 14365 52144 14399
rect 52092 14356 52144 14365
rect 52276 14399 52328 14408
rect 52276 14365 52285 14399
rect 52285 14365 52319 14399
rect 52319 14365 52328 14399
rect 52276 14356 52328 14365
rect 52460 14356 52512 14408
rect 52736 14356 52788 14408
rect 46296 14220 46348 14272
rect 48320 14288 48372 14340
rect 49056 14220 49108 14272
rect 51540 14288 51592 14340
rect 53288 14399 53340 14408
rect 53288 14365 53297 14399
rect 53297 14365 53331 14399
rect 53331 14365 53340 14399
rect 53288 14356 53340 14365
rect 53840 14356 53892 14408
rect 54576 14356 54628 14408
rect 55680 14399 55732 14408
rect 55680 14365 55689 14399
rect 55689 14365 55723 14399
rect 55723 14365 55732 14399
rect 55680 14356 55732 14365
rect 57888 14356 57940 14408
rect 50344 14220 50396 14272
rect 52276 14220 52328 14272
rect 53104 14220 53156 14272
rect 54392 14220 54444 14272
rect 54852 14263 54904 14272
rect 54852 14229 54861 14263
rect 54861 14229 54895 14263
rect 54895 14229 54904 14263
rect 54852 14220 54904 14229
rect 56692 14263 56744 14272
rect 56692 14229 56701 14263
rect 56701 14229 56735 14263
rect 56735 14229 56744 14263
rect 56692 14220 56744 14229
rect 57796 14263 57848 14272
rect 57796 14229 57805 14263
rect 57805 14229 57839 14263
rect 57839 14229 57848 14263
rect 57796 14220 57848 14229
rect 58072 14220 58124 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 28724 14059 28776 14068
rect 26424 13948 26476 14000
rect 27896 13948 27948 14000
rect 24952 13923 25004 13932
rect 24952 13889 24961 13923
rect 24961 13889 24995 13923
rect 24995 13889 25004 13923
rect 24952 13880 25004 13889
rect 25780 13880 25832 13932
rect 26148 13880 26200 13932
rect 26516 13880 26568 13932
rect 26976 13880 27028 13932
rect 28724 14025 28733 14059
rect 28733 14025 28767 14059
rect 28767 14025 28776 14059
rect 28724 14016 28776 14025
rect 30012 14016 30064 14068
rect 30380 14016 30432 14068
rect 28816 13923 28868 13932
rect 25964 13744 26016 13796
rect 26240 13812 26292 13864
rect 26884 13744 26936 13796
rect 26056 13676 26108 13728
rect 28816 13889 28825 13923
rect 28825 13889 28859 13923
rect 28859 13889 28868 13923
rect 28816 13880 28868 13889
rect 29368 13923 29420 13932
rect 29368 13889 29377 13923
rect 29377 13889 29411 13923
rect 29411 13889 29420 13923
rect 29368 13880 29420 13889
rect 29552 13923 29604 13932
rect 29552 13889 29561 13923
rect 29561 13889 29595 13923
rect 29595 13889 29604 13923
rect 29552 13880 29604 13889
rect 29736 13948 29788 14000
rect 31300 14016 31352 14068
rect 32496 14016 32548 14068
rect 33600 14016 33652 14068
rect 33692 14016 33744 14068
rect 35716 14016 35768 14068
rect 29920 13923 29972 13932
rect 29920 13889 29929 13923
rect 29929 13889 29963 13923
rect 29963 13889 29972 13923
rect 29920 13880 29972 13889
rect 31024 13923 31076 13932
rect 31024 13889 31033 13923
rect 31033 13889 31067 13923
rect 31067 13889 31076 13923
rect 31024 13880 31076 13889
rect 31668 13880 31720 13932
rect 32588 13880 32640 13932
rect 32956 13880 33008 13932
rect 33416 13923 33468 13932
rect 33416 13889 33425 13923
rect 33425 13889 33459 13923
rect 33459 13889 33468 13923
rect 33416 13880 33468 13889
rect 28724 13812 28776 13864
rect 31760 13812 31812 13864
rect 32220 13812 32272 13864
rect 33324 13855 33376 13864
rect 33324 13821 33333 13855
rect 33333 13821 33367 13855
rect 33367 13821 33376 13855
rect 33324 13812 33376 13821
rect 33876 13880 33928 13932
rect 37004 14016 37056 14068
rect 37280 14016 37332 14068
rect 38660 14016 38712 14068
rect 38844 14016 38896 14068
rect 41604 14059 41656 14068
rect 41604 14025 41613 14059
rect 41613 14025 41647 14059
rect 41647 14025 41656 14059
rect 41604 14016 41656 14025
rect 43536 14016 43588 14068
rect 37372 13948 37424 14000
rect 38476 13948 38528 14000
rect 34520 13880 34572 13932
rect 34704 13923 34756 13932
rect 34704 13889 34713 13923
rect 34713 13889 34747 13923
rect 34747 13889 34756 13923
rect 34704 13880 34756 13889
rect 35440 13880 35492 13932
rect 35808 13923 35860 13932
rect 35808 13889 35817 13923
rect 35817 13889 35851 13923
rect 35851 13889 35860 13923
rect 35808 13880 35860 13889
rect 36084 13812 36136 13864
rect 36268 13880 36320 13932
rect 36912 13923 36964 13932
rect 36360 13812 36412 13864
rect 28908 13744 28960 13796
rect 29460 13676 29512 13728
rect 33508 13744 33560 13796
rect 36912 13889 36921 13923
rect 36921 13889 36955 13923
rect 36955 13889 36964 13923
rect 36912 13880 36964 13889
rect 39212 13923 39264 13932
rect 37188 13812 37240 13864
rect 39212 13889 39221 13923
rect 39221 13889 39255 13923
rect 39255 13889 39264 13923
rect 39212 13880 39264 13889
rect 39856 13923 39908 13932
rect 39856 13889 39865 13923
rect 39865 13889 39899 13923
rect 39899 13889 39908 13923
rect 39856 13880 39908 13889
rect 42984 13948 43036 14000
rect 40500 13923 40552 13932
rect 40500 13889 40509 13923
rect 40509 13889 40543 13923
rect 40543 13889 40552 13923
rect 40500 13880 40552 13889
rect 39120 13812 39172 13864
rect 40408 13812 40460 13864
rect 43352 13880 43404 13932
rect 41696 13812 41748 13864
rect 42340 13812 42392 13864
rect 44364 13880 44416 13932
rect 44548 13880 44600 13932
rect 45284 13880 45336 13932
rect 45376 13923 45428 13932
rect 45376 13889 45385 13923
rect 45385 13889 45419 13923
rect 45419 13889 45428 13923
rect 45376 13880 45428 13889
rect 44824 13812 44876 13864
rect 45928 14016 45980 14068
rect 46848 14016 46900 14068
rect 47032 14016 47084 14068
rect 47400 14016 47452 14068
rect 47860 14016 47912 14068
rect 45836 13880 45888 13932
rect 46204 13880 46256 13932
rect 50160 13948 50212 14000
rect 52092 14016 52144 14068
rect 52368 14016 52420 14068
rect 53380 14016 53432 14068
rect 54668 14016 54720 14068
rect 55128 14059 55180 14068
rect 55128 14025 55137 14059
rect 55137 14025 55171 14059
rect 55171 14025 55180 14059
rect 55128 14016 55180 14025
rect 55220 14016 55272 14068
rect 46664 13923 46716 13932
rect 38476 13744 38528 13796
rect 43536 13744 43588 13796
rect 31116 13676 31168 13728
rect 32128 13676 32180 13728
rect 37924 13676 37976 13728
rect 39212 13676 39264 13728
rect 40224 13676 40276 13728
rect 44640 13719 44692 13728
rect 44640 13685 44649 13719
rect 44649 13685 44683 13719
rect 44683 13685 44692 13719
rect 44640 13676 44692 13685
rect 46664 13889 46673 13923
rect 46673 13889 46707 13923
rect 46707 13889 46716 13923
rect 46664 13880 46716 13889
rect 46848 13923 46900 13932
rect 46848 13889 46857 13923
rect 46857 13889 46891 13923
rect 46891 13889 46900 13923
rect 46848 13880 46900 13889
rect 47400 13880 47452 13932
rect 48504 13880 48556 13932
rect 46756 13855 46808 13864
rect 46756 13821 46765 13855
rect 46765 13821 46799 13855
rect 46799 13821 46808 13855
rect 46756 13812 46808 13821
rect 47768 13855 47820 13864
rect 47768 13821 47777 13855
rect 47777 13821 47811 13855
rect 47811 13821 47820 13855
rect 47768 13812 47820 13821
rect 49424 13812 49476 13864
rect 49976 13812 50028 13864
rect 50160 13855 50212 13864
rect 50160 13821 50169 13855
rect 50169 13821 50203 13855
rect 50203 13821 50212 13855
rect 50160 13812 50212 13821
rect 51540 13948 51592 14000
rect 54852 13948 54904 14000
rect 55496 13948 55548 14000
rect 50620 13880 50672 13932
rect 51264 13923 51316 13932
rect 51264 13889 51273 13923
rect 51273 13889 51307 13923
rect 51307 13889 51316 13923
rect 51264 13880 51316 13889
rect 51632 13880 51684 13932
rect 52276 13880 52328 13932
rect 49056 13744 49108 13796
rect 50436 13855 50488 13864
rect 50436 13821 50445 13855
rect 50445 13821 50479 13855
rect 50479 13821 50488 13855
rect 50436 13812 50488 13821
rect 52828 13812 52880 13864
rect 51172 13744 51224 13796
rect 52184 13744 52236 13796
rect 54208 13923 54260 13932
rect 54208 13889 54217 13923
rect 54217 13889 54251 13923
rect 54251 13889 54260 13923
rect 54208 13880 54260 13889
rect 54576 13923 54628 13932
rect 54576 13889 54585 13923
rect 54585 13889 54619 13923
rect 54619 13889 54628 13923
rect 54576 13880 54628 13889
rect 56232 14016 56284 14068
rect 57612 14016 57664 14068
rect 58072 14059 58124 14068
rect 58072 14025 58081 14059
rect 58081 14025 58115 14059
rect 58115 14025 58124 14059
rect 58072 14016 58124 14025
rect 56048 13923 56100 13932
rect 56048 13889 56057 13923
rect 56057 13889 56091 13923
rect 56091 13889 56100 13923
rect 56048 13880 56100 13889
rect 56416 13880 56468 13932
rect 57336 13948 57388 14000
rect 53288 13812 53340 13864
rect 53932 13812 53984 13864
rect 56508 13812 56560 13864
rect 53380 13744 53432 13796
rect 57796 13744 57848 13796
rect 48412 13676 48464 13728
rect 48964 13676 49016 13728
rect 49608 13676 49660 13728
rect 52920 13676 52972 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 24952 13515 25004 13524
rect 24952 13481 24961 13515
rect 24961 13481 24995 13515
rect 24995 13481 25004 13515
rect 24952 13472 25004 13481
rect 25688 13515 25740 13524
rect 25688 13481 25697 13515
rect 25697 13481 25731 13515
rect 25731 13481 25740 13515
rect 25688 13472 25740 13481
rect 26240 13472 26292 13524
rect 31300 13515 31352 13524
rect 26884 13404 26936 13456
rect 27804 13404 27856 13456
rect 26056 13336 26108 13388
rect 31300 13481 31309 13515
rect 31309 13481 31343 13515
rect 31343 13481 31352 13515
rect 31300 13472 31352 13481
rect 32128 13472 32180 13524
rect 33876 13472 33928 13524
rect 36728 13472 36780 13524
rect 37188 13472 37240 13524
rect 37372 13472 37424 13524
rect 38108 13472 38160 13524
rect 39212 13515 39264 13524
rect 39212 13481 39221 13515
rect 39221 13481 39255 13515
rect 39255 13481 39264 13515
rect 39212 13472 39264 13481
rect 40316 13472 40368 13524
rect 43076 13515 43128 13524
rect 43076 13481 43085 13515
rect 43085 13481 43119 13515
rect 43119 13481 43128 13515
rect 43076 13472 43128 13481
rect 44272 13515 44324 13524
rect 44272 13481 44281 13515
rect 44281 13481 44315 13515
rect 44315 13481 44324 13515
rect 46388 13515 46440 13524
rect 44272 13472 44324 13481
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 25964 13268 26016 13320
rect 26884 13311 26936 13320
rect 26884 13277 26893 13311
rect 26893 13277 26927 13311
rect 26927 13277 26936 13311
rect 26884 13268 26936 13277
rect 27804 13311 27856 13320
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 29092 13336 29144 13388
rect 31668 13404 31720 13456
rect 33600 13404 33652 13456
rect 39120 13404 39172 13456
rect 28908 13311 28960 13320
rect 24860 13243 24912 13252
rect 24860 13209 24869 13243
rect 24869 13209 24903 13243
rect 24903 13209 24912 13243
rect 24860 13200 24912 13209
rect 26976 13243 27028 13252
rect 26976 13209 26985 13243
rect 26985 13209 27019 13243
rect 27019 13209 27028 13243
rect 26976 13200 27028 13209
rect 24492 13132 24544 13184
rect 27712 13132 27764 13184
rect 28908 13277 28917 13311
rect 28917 13277 28951 13311
rect 28951 13277 28960 13311
rect 28908 13268 28960 13277
rect 29000 13311 29052 13320
rect 29000 13277 29009 13311
rect 29009 13277 29043 13311
rect 29043 13277 29052 13311
rect 29000 13268 29052 13277
rect 29368 13268 29420 13320
rect 29828 13268 29880 13320
rect 30840 13311 30892 13320
rect 30840 13277 30849 13311
rect 30849 13277 30883 13311
rect 30883 13277 30892 13311
rect 30840 13268 30892 13277
rect 33048 13336 33100 13388
rect 33232 13311 33284 13320
rect 30748 13200 30800 13252
rect 33232 13277 33241 13311
rect 33241 13277 33275 13311
rect 33275 13277 33284 13311
rect 33232 13268 33284 13277
rect 33968 13268 34020 13320
rect 34244 13311 34296 13320
rect 34244 13277 34253 13311
rect 34253 13277 34287 13311
rect 34287 13277 34296 13311
rect 34244 13268 34296 13277
rect 35164 13200 35216 13252
rect 29184 13132 29236 13184
rect 33508 13132 33560 13184
rect 34336 13132 34388 13184
rect 37188 13336 37240 13388
rect 38660 13336 38712 13388
rect 40408 13336 40460 13388
rect 41236 13336 41288 13388
rect 43352 13336 43404 13388
rect 35440 13311 35492 13320
rect 35440 13277 35449 13311
rect 35449 13277 35483 13311
rect 35483 13277 35492 13311
rect 35440 13268 35492 13277
rect 36176 13268 36228 13320
rect 41972 13311 42024 13320
rect 36728 13200 36780 13252
rect 36820 13200 36872 13252
rect 41972 13277 41981 13311
rect 41981 13277 42015 13311
rect 42015 13277 42024 13311
rect 41972 13268 42024 13277
rect 42984 13311 43036 13320
rect 40224 13200 40276 13252
rect 42984 13277 42993 13311
rect 42993 13277 43027 13311
rect 43027 13277 43036 13311
rect 42984 13268 43036 13277
rect 43168 13311 43220 13320
rect 43168 13277 43177 13311
rect 43177 13277 43211 13311
rect 43211 13277 43220 13311
rect 43168 13268 43220 13277
rect 44364 13404 44416 13456
rect 45928 13404 45980 13456
rect 46020 13404 46072 13456
rect 46388 13481 46397 13515
rect 46397 13481 46431 13515
rect 46431 13481 46440 13515
rect 46388 13472 46440 13481
rect 47124 13472 47176 13524
rect 48044 13472 48096 13524
rect 48504 13472 48556 13524
rect 48688 13515 48740 13524
rect 48688 13481 48697 13515
rect 48697 13481 48731 13515
rect 48731 13481 48740 13515
rect 48688 13472 48740 13481
rect 47216 13404 47268 13456
rect 50068 13472 50120 13524
rect 50436 13472 50488 13524
rect 50988 13472 51040 13524
rect 51356 13472 51408 13524
rect 52184 13515 52236 13524
rect 52184 13481 52193 13515
rect 52193 13481 52227 13515
rect 52227 13481 52236 13515
rect 52184 13472 52236 13481
rect 52828 13472 52880 13524
rect 54392 13472 54444 13524
rect 54576 13472 54628 13524
rect 43904 13336 43956 13388
rect 43812 13311 43864 13320
rect 43812 13277 43819 13311
rect 43819 13277 43864 13311
rect 43812 13268 43864 13277
rect 44548 13336 44600 13388
rect 44640 13268 44692 13320
rect 45376 13268 45428 13320
rect 46388 13336 46440 13388
rect 46756 13336 46808 13388
rect 48964 13404 49016 13456
rect 47952 13336 48004 13388
rect 48504 13336 48556 13388
rect 38016 13132 38068 13184
rect 38292 13132 38344 13184
rect 38568 13132 38620 13184
rect 40776 13132 40828 13184
rect 42340 13175 42392 13184
rect 42340 13141 42349 13175
rect 42349 13141 42383 13175
rect 42383 13141 42392 13175
rect 42340 13132 42392 13141
rect 45652 13200 45704 13252
rect 45192 13175 45244 13184
rect 45192 13141 45201 13175
rect 45201 13141 45235 13175
rect 45235 13141 45244 13175
rect 45192 13132 45244 13141
rect 47032 13200 47084 13252
rect 48136 13268 48188 13320
rect 48228 13268 48280 13320
rect 54208 13404 54260 13456
rect 49700 13336 49752 13388
rect 48044 13200 48096 13252
rect 46204 13132 46256 13184
rect 48504 13243 48556 13252
rect 48504 13209 48513 13243
rect 48513 13209 48547 13243
rect 48547 13209 48556 13243
rect 48504 13200 48556 13209
rect 48688 13200 48740 13252
rect 49792 13268 49844 13320
rect 51356 13336 51408 13388
rect 50712 13268 50764 13320
rect 51816 13336 51868 13388
rect 52644 13336 52696 13388
rect 53748 13336 53800 13388
rect 49700 13200 49752 13252
rect 52460 13268 52512 13320
rect 53196 13268 53248 13320
rect 53472 13268 53524 13320
rect 55128 13404 55180 13456
rect 55588 13404 55640 13456
rect 56508 13472 56560 13524
rect 56600 13515 56652 13524
rect 56600 13481 56609 13515
rect 56609 13481 56643 13515
rect 56643 13481 56652 13515
rect 56600 13472 56652 13481
rect 56416 13404 56468 13456
rect 56232 13268 56284 13320
rect 57980 13268 58032 13320
rect 58440 13268 58492 13320
rect 49608 13132 49660 13184
rect 51172 13132 51224 13184
rect 51448 13132 51500 13184
rect 52552 13132 52604 13184
rect 53196 13132 53248 13184
rect 53656 13132 53708 13184
rect 54208 13243 54260 13252
rect 54208 13209 54217 13243
rect 54217 13209 54251 13243
rect 54251 13209 54260 13243
rect 54208 13200 54260 13209
rect 56048 13200 56100 13252
rect 55864 13132 55916 13184
rect 56232 13132 56284 13184
rect 58256 13175 58308 13184
rect 58256 13141 58265 13175
rect 58265 13141 58299 13175
rect 58299 13141 58308 13175
rect 58256 13132 58308 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 25872 12971 25924 12980
rect 25872 12937 25881 12971
rect 25881 12937 25915 12971
rect 25915 12937 25924 12971
rect 25872 12928 25924 12937
rect 26148 12928 26200 12980
rect 27896 12928 27948 12980
rect 28908 12928 28960 12980
rect 29184 12928 29236 12980
rect 31852 12928 31904 12980
rect 33416 12928 33468 12980
rect 34244 12971 34296 12980
rect 34244 12937 34253 12971
rect 34253 12937 34287 12971
rect 34287 12937 34296 12971
rect 34244 12928 34296 12937
rect 34520 12928 34572 12980
rect 35348 12928 35400 12980
rect 35900 12928 35952 12980
rect 36452 12928 36504 12980
rect 37924 12928 37976 12980
rect 40224 12928 40276 12980
rect 40500 12928 40552 12980
rect 42708 12971 42760 12980
rect 42708 12937 42717 12971
rect 42717 12937 42751 12971
rect 42751 12937 42760 12971
rect 42708 12928 42760 12937
rect 1860 12588 1912 12640
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 24860 12792 24912 12844
rect 24492 12724 24544 12776
rect 25964 12792 26016 12844
rect 26056 12835 26108 12844
rect 26056 12801 26065 12835
rect 26065 12801 26099 12835
rect 26099 12801 26108 12835
rect 26056 12792 26108 12801
rect 26424 12792 26476 12844
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 27436 12835 27488 12844
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 27712 12835 27764 12844
rect 27712 12801 27721 12835
rect 27721 12801 27755 12835
rect 27755 12801 27764 12835
rect 27712 12792 27764 12801
rect 28080 12860 28132 12912
rect 28172 12792 28224 12844
rect 29092 12792 29144 12844
rect 29460 12792 29512 12844
rect 29828 12835 29880 12844
rect 29828 12801 29837 12835
rect 29837 12801 29871 12835
rect 29871 12801 29880 12835
rect 29828 12792 29880 12801
rect 30104 12792 30156 12844
rect 27988 12724 28040 12776
rect 27252 12656 27304 12708
rect 27344 12656 27396 12708
rect 29552 12724 29604 12776
rect 32496 12767 32548 12776
rect 32496 12733 32505 12767
rect 32505 12733 32539 12767
rect 32539 12733 32548 12767
rect 32496 12724 32548 12733
rect 32588 12767 32640 12776
rect 32588 12733 32597 12767
rect 32597 12733 32631 12767
rect 32631 12733 32640 12767
rect 32588 12724 32640 12733
rect 33600 12835 33652 12844
rect 33600 12801 33609 12835
rect 33609 12801 33643 12835
rect 33643 12801 33652 12835
rect 33600 12792 33652 12801
rect 33968 12792 34020 12844
rect 34336 12792 34388 12844
rect 34980 12835 35032 12844
rect 34980 12801 34989 12835
rect 34989 12801 35023 12835
rect 35023 12801 35032 12835
rect 34980 12792 35032 12801
rect 35164 12835 35216 12844
rect 35164 12801 35173 12835
rect 35173 12801 35207 12835
rect 35207 12801 35216 12835
rect 35164 12792 35216 12801
rect 35716 12792 35768 12844
rect 32864 12656 32916 12708
rect 35348 12767 35400 12776
rect 35348 12733 35357 12767
rect 35357 12733 35391 12767
rect 35391 12733 35400 12767
rect 35900 12792 35952 12844
rect 36084 12792 36136 12844
rect 36268 12792 36320 12844
rect 36544 12835 36596 12844
rect 36544 12801 36553 12835
rect 36553 12801 36587 12835
rect 36587 12801 36596 12835
rect 36544 12792 36596 12801
rect 36636 12835 36688 12844
rect 36636 12801 36645 12835
rect 36645 12801 36679 12835
rect 36679 12801 36688 12835
rect 36636 12792 36688 12801
rect 37188 12792 37240 12844
rect 39396 12860 39448 12912
rect 42616 12860 42668 12912
rect 44548 12928 44600 12980
rect 44916 12928 44968 12980
rect 45928 12928 45980 12980
rect 47308 12928 47360 12980
rect 43904 12860 43956 12912
rect 44640 12860 44692 12912
rect 46020 12860 46072 12912
rect 48228 12860 48280 12912
rect 48412 12860 48464 12912
rect 49608 12928 49660 12980
rect 49884 12928 49936 12980
rect 38292 12792 38344 12844
rect 35348 12724 35400 12733
rect 26792 12588 26844 12640
rect 28724 12588 28776 12640
rect 30380 12588 30432 12640
rect 30748 12588 30800 12640
rect 31024 12588 31076 12640
rect 34152 12588 34204 12640
rect 36084 12656 36136 12708
rect 37004 12724 37056 12776
rect 38936 12767 38988 12776
rect 38936 12733 38945 12767
rect 38945 12733 38979 12767
rect 38979 12733 38988 12767
rect 38936 12724 38988 12733
rect 39212 12792 39264 12844
rect 42892 12835 42944 12844
rect 40684 12724 40736 12776
rect 42892 12801 42901 12835
rect 42901 12801 42935 12835
rect 42935 12801 42944 12835
rect 42892 12792 42944 12801
rect 43076 12792 43128 12844
rect 43260 12792 43312 12844
rect 43628 12792 43680 12844
rect 45376 12792 45428 12844
rect 47216 12792 47268 12844
rect 48044 12835 48096 12844
rect 48044 12801 48053 12835
rect 48053 12801 48087 12835
rect 48087 12801 48096 12835
rect 48044 12792 48096 12801
rect 48320 12792 48372 12844
rect 49792 12860 49844 12912
rect 53840 12928 53892 12980
rect 41972 12724 42024 12776
rect 45192 12724 45244 12776
rect 46664 12724 46716 12776
rect 46756 12767 46808 12776
rect 46756 12733 46765 12767
rect 46765 12733 46799 12767
rect 46799 12733 46808 12767
rect 49240 12801 49249 12806
rect 49249 12801 49283 12806
rect 49283 12801 49292 12806
rect 49240 12754 49292 12801
rect 49424 12835 49476 12844
rect 49424 12801 49438 12835
rect 49438 12801 49472 12835
rect 49472 12801 49476 12835
rect 52092 12860 52144 12912
rect 52552 12860 52604 12912
rect 50620 12835 50672 12844
rect 49424 12792 49476 12801
rect 50620 12801 50629 12835
rect 50629 12801 50663 12835
rect 50663 12801 50672 12835
rect 50620 12792 50672 12801
rect 51908 12792 51960 12844
rect 46756 12724 46808 12733
rect 40132 12656 40184 12708
rect 40408 12656 40460 12708
rect 44548 12699 44600 12708
rect 44548 12665 44557 12699
rect 44557 12665 44591 12699
rect 44591 12665 44600 12699
rect 44548 12656 44600 12665
rect 44640 12656 44692 12708
rect 44916 12656 44968 12708
rect 37188 12588 37240 12640
rect 39304 12588 39356 12640
rect 40040 12631 40092 12640
rect 40040 12597 40049 12631
rect 40049 12597 40083 12631
rect 40083 12597 40092 12631
rect 40040 12588 40092 12597
rect 43720 12588 43772 12640
rect 46388 12588 46440 12640
rect 46664 12588 46716 12640
rect 48136 12588 48188 12640
rect 49792 12724 49844 12776
rect 50988 12724 51040 12776
rect 51356 12724 51408 12776
rect 52460 12792 52512 12844
rect 52920 12835 52972 12844
rect 52920 12801 52929 12835
rect 52929 12801 52963 12835
rect 52963 12801 52972 12835
rect 52920 12792 52972 12801
rect 53104 12792 53156 12844
rect 56232 12860 56284 12912
rect 56968 12860 57020 12912
rect 57888 12860 57940 12912
rect 54852 12835 54904 12844
rect 53748 12724 53800 12776
rect 54852 12801 54861 12835
rect 54861 12801 54895 12835
rect 54895 12801 54904 12835
rect 54852 12792 54904 12801
rect 55036 12835 55088 12844
rect 55036 12801 55045 12835
rect 55045 12801 55079 12835
rect 55079 12801 55088 12835
rect 55036 12792 55088 12801
rect 54944 12724 54996 12776
rect 55772 12767 55824 12776
rect 55772 12733 55781 12767
rect 55781 12733 55815 12767
rect 55815 12733 55824 12767
rect 55772 12724 55824 12733
rect 49976 12656 50028 12708
rect 51080 12656 51132 12708
rect 52092 12656 52144 12708
rect 54392 12656 54444 12708
rect 49608 12631 49660 12640
rect 49608 12597 49617 12631
rect 49617 12597 49651 12631
rect 49651 12597 49660 12631
rect 49608 12588 49660 12597
rect 53564 12588 53616 12640
rect 55404 12588 55456 12640
rect 55680 12631 55732 12640
rect 55680 12597 55689 12631
rect 55689 12597 55723 12631
rect 55723 12597 55732 12631
rect 56968 12656 57020 12708
rect 55680 12588 55732 12597
rect 56692 12588 56744 12640
rect 57428 12631 57480 12640
rect 57428 12597 57437 12631
rect 57437 12597 57471 12631
rect 57471 12597 57480 12631
rect 57428 12588 57480 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 24492 12384 24544 12436
rect 25780 12384 25832 12436
rect 27436 12384 27488 12436
rect 25688 12316 25740 12368
rect 27344 12291 27396 12300
rect 27344 12257 27353 12291
rect 27353 12257 27387 12291
rect 27387 12257 27396 12291
rect 27344 12248 27396 12257
rect 27436 12291 27488 12300
rect 27436 12257 27445 12291
rect 27445 12257 27479 12291
rect 27479 12257 27488 12291
rect 28816 12316 28868 12368
rect 30380 12316 30432 12368
rect 32496 12384 32548 12436
rect 33140 12427 33192 12436
rect 33140 12393 33149 12427
rect 33149 12393 33183 12427
rect 33183 12393 33192 12427
rect 33140 12384 33192 12393
rect 36636 12384 36688 12436
rect 37188 12384 37240 12436
rect 32404 12316 32456 12368
rect 27436 12248 27488 12257
rect 27528 12223 27580 12232
rect 27528 12189 27537 12223
rect 27537 12189 27571 12223
rect 27571 12189 27580 12223
rect 27528 12180 27580 12189
rect 28724 12223 28776 12232
rect 28724 12189 28733 12223
rect 28733 12189 28767 12223
rect 28767 12189 28776 12223
rect 28724 12180 28776 12189
rect 33324 12291 33376 12300
rect 33324 12257 33333 12291
rect 33333 12257 33367 12291
rect 33367 12257 33376 12291
rect 33324 12248 33376 12257
rect 26792 12112 26844 12164
rect 28080 12112 28132 12164
rect 28356 12112 28408 12164
rect 26608 12087 26660 12096
rect 26608 12053 26617 12087
rect 26617 12053 26651 12087
rect 26651 12053 26660 12087
rect 26608 12044 26660 12053
rect 26884 12044 26936 12096
rect 28632 12044 28684 12096
rect 30196 12180 30248 12232
rect 30288 12223 30340 12232
rect 30288 12189 30297 12223
rect 30297 12189 30331 12223
rect 30331 12189 30340 12223
rect 30288 12180 30340 12189
rect 30012 12112 30064 12164
rect 30380 12112 30432 12164
rect 30748 12180 30800 12232
rect 33048 12180 33100 12232
rect 33416 12223 33468 12232
rect 33416 12189 33425 12223
rect 33425 12189 33459 12223
rect 33459 12189 33468 12223
rect 33416 12180 33468 12189
rect 31852 12112 31904 12164
rect 34428 12248 34480 12300
rect 33692 12223 33744 12232
rect 33692 12189 33701 12223
rect 33701 12189 33735 12223
rect 33735 12189 33744 12223
rect 33692 12180 33744 12189
rect 33876 12180 33928 12232
rect 35072 12180 35124 12232
rect 37740 12248 37792 12300
rect 38844 12384 38896 12436
rect 39396 12384 39448 12436
rect 40592 12427 40644 12436
rect 37924 12316 37976 12368
rect 36360 12180 36412 12232
rect 36728 12180 36780 12232
rect 37648 12223 37700 12232
rect 29276 12044 29328 12096
rect 30748 12044 30800 12096
rect 31944 12044 31996 12096
rect 33784 12155 33836 12164
rect 33784 12121 33793 12155
rect 33793 12121 33827 12155
rect 33827 12121 33836 12155
rect 33784 12112 33836 12121
rect 34060 12112 34112 12164
rect 37280 12112 37332 12164
rect 37648 12189 37657 12223
rect 37657 12189 37691 12223
rect 37691 12189 37700 12223
rect 37648 12180 37700 12189
rect 37924 12223 37976 12232
rect 37924 12189 37933 12223
rect 37933 12189 37967 12223
rect 37967 12189 37976 12223
rect 37924 12180 37976 12189
rect 38108 12180 38160 12232
rect 40040 12316 40092 12368
rect 40592 12393 40601 12427
rect 40601 12393 40635 12427
rect 40635 12393 40644 12427
rect 40592 12384 40644 12393
rect 44088 12384 44140 12436
rect 46112 12384 46164 12436
rect 48136 12384 48188 12436
rect 48596 12384 48648 12436
rect 48780 12384 48832 12436
rect 50712 12384 50764 12436
rect 52092 12384 52144 12436
rect 53656 12384 53708 12436
rect 54024 12384 54076 12436
rect 54944 12384 54996 12436
rect 58072 12384 58124 12436
rect 40684 12316 40736 12368
rect 43168 12316 43220 12368
rect 43720 12316 43772 12368
rect 44916 12316 44968 12368
rect 45284 12316 45336 12368
rect 48320 12316 48372 12368
rect 40132 12223 40184 12232
rect 40132 12189 40141 12223
rect 40141 12189 40175 12223
rect 40175 12189 40184 12223
rect 40132 12180 40184 12189
rect 40316 12223 40368 12232
rect 40316 12189 40325 12223
rect 40325 12189 40359 12223
rect 40359 12189 40368 12223
rect 40316 12180 40368 12189
rect 40408 12223 40460 12232
rect 40408 12189 40417 12223
rect 40417 12189 40451 12223
rect 40451 12189 40460 12223
rect 43536 12248 43588 12300
rect 45560 12248 45612 12300
rect 45928 12248 45980 12300
rect 40408 12180 40460 12189
rect 43168 12223 43220 12232
rect 43168 12189 43177 12223
rect 43177 12189 43211 12223
rect 43211 12189 43220 12223
rect 43168 12180 43220 12189
rect 43076 12112 43128 12164
rect 43352 12223 43404 12232
rect 43352 12189 43361 12223
rect 43361 12189 43395 12223
rect 43395 12189 43404 12223
rect 43352 12180 43404 12189
rect 45468 12223 45520 12232
rect 45468 12189 45477 12223
rect 45477 12189 45511 12223
rect 45511 12189 45520 12223
rect 48136 12248 48188 12300
rect 48504 12316 48556 12368
rect 49424 12316 49476 12368
rect 45468 12180 45520 12189
rect 43996 12112 44048 12164
rect 45284 12112 45336 12164
rect 45652 12112 45704 12164
rect 46112 12112 46164 12164
rect 46296 12112 46348 12164
rect 32404 12044 32456 12096
rect 34888 12044 34940 12096
rect 35256 12044 35308 12096
rect 35900 12044 35952 12096
rect 36176 12044 36228 12096
rect 36636 12044 36688 12096
rect 36820 12044 36872 12096
rect 37648 12044 37700 12096
rect 38108 12044 38160 12096
rect 38568 12044 38620 12096
rect 40960 12044 41012 12096
rect 41236 12044 41288 12096
rect 43260 12044 43312 12096
rect 44180 12087 44232 12096
rect 44180 12053 44189 12087
rect 44189 12053 44223 12087
rect 44223 12053 44232 12087
rect 44180 12044 44232 12053
rect 45468 12044 45520 12096
rect 45560 12044 45612 12096
rect 47032 12223 47084 12232
rect 47032 12189 47041 12223
rect 47041 12189 47075 12223
rect 47075 12189 47084 12223
rect 47032 12180 47084 12189
rect 48964 12248 49016 12300
rect 46664 12155 46716 12164
rect 46664 12121 46673 12155
rect 46673 12121 46707 12155
rect 46707 12121 46716 12155
rect 46664 12112 46716 12121
rect 46848 12155 46900 12164
rect 46848 12121 46883 12155
rect 46883 12121 46900 12155
rect 46848 12112 46900 12121
rect 47124 12112 47176 12164
rect 48596 12223 48648 12232
rect 48596 12189 48605 12223
rect 48605 12189 48639 12223
rect 48639 12189 48648 12223
rect 49700 12248 49752 12300
rect 50344 12248 50396 12300
rect 52736 12316 52788 12368
rect 53380 12359 53432 12368
rect 53380 12325 53389 12359
rect 53389 12325 53423 12359
rect 53423 12325 53432 12359
rect 53380 12316 53432 12325
rect 54484 12316 54536 12368
rect 55496 12359 55548 12368
rect 55496 12325 55505 12359
rect 55505 12325 55539 12359
rect 55539 12325 55548 12359
rect 55496 12316 55548 12325
rect 48596 12180 48648 12189
rect 48964 12112 49016 12164
rect 49608 12223 49660 12232
rect 49608 12189 49617 12223
rect 49617 12189 49651 12223
rect 49651 12189 49660 12223
rect 49608 12180 49660 12189
rect 49976 12180 50028 12232
rect 50436 12112 50488 12164
rect 52184 12180 52236 12232
rect 51632 12112 51684 12164
rect 52368 12180 52420 12232
rect 52552 12223 52604 12232
rect 52552 12189 52561 12223
rect 52561 12189 52595 12223
rect 52595 12189 52604 12223
rect 53288 12248 53340 12300
rect 53656 12248 53708 12300
rect 55956 12248 56008 12300
rect 52552 12180 52604 12189
rect 52828 12180 52880 12232
rect 53564 12223 53616 12232
rect 53564 12189 53573 12223
rect 53573 12189 53607 12223
rect 53607 12189 53616 12223
rect 53564 12180 53616 12189
rect 53840 12180 53892 12232
rect 54668 12180 54720 12232
rect 52920 12112 52972 12164
rect 55220 12180 55272 12232
rect 55680 12180 55732 12232
rect 55496 12112 55548 12164
rect 48228 12044 48280 12096
rect 48596 12044 48648 12096
rect 49424 12044 49476 12096
rect 50804 12044 50856 12096
rect 53564 12044 53616 12096
rect 54208 12044 54260 12096
rect 54852 12044 54904 12096
rect 55312 12044 55364 12096
rect 55680 12044 55732 12096
rect 57336 12087 57388 12096
rect 57336 12053 57345 12087
rect 57345 12053 57379 12087
rect 57379 12053 57388 12087
rect 57336 12044 57388 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 24768 11883 24820 11892
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 24952 11840 25004 11892
rect 24032 11772 24084 11824
rect 1676 11611 1728 11620
rect 1676 11577 1685 11611
rect 1685 11577 1719 11611
rect 1719 11577 1728 11611
rect 1676 11568 1728 11577
rect 24952 11704 25004 11756
rect 25228 11772 25280 11824
rect 27896 11840 27948 11892
rect 29184 11883 29236 11892
rect 29184 11849 29193 11883
rect 29193 11849 29227 11883
rect 29227 11849 29236 11883
rect 29184 11840 29236 11849
rect 33416 11840 33468 11892
rect 33784 11840 33836 11892
rect 34060 11840 34112 11892
rect 27160 11815 27212 11824
rect 27160 11781 27169 11815
rect 27169 11781 27203 11815
rect 27203 11781 27212 11815
rect 27160 11772 27212 11781
rect 28080 11772 28132 11824
rect 31024 11815 31076 11824
rect 31024 11781 31033 11815
rect 31033 11781 31067 11815
rect 31067 11781 31076 11815
rect 31024 11772 31076 11781
rect 31852 11772 31904 11824
rect 33876 11815 33928 11824
rect 33876 11781 33885 11815
rect 33885 11781 33919 11815
rect 33919 11781 33928 11815
rect 33876 11772 33928 11781
rect 35808 11840 35860 11892
rect 25688 11747 25740 11756
rect 24400 11568 24452 11620
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 26056 11747 26108 11756
rect 26056 11713 26065 11747
rect 26065 11713 26099 11747
rect 26099 11713 26108 11747
rect 26056 11704 26108 11713
rect 27436 11704 27488 11756
rect 28264 11704 28316 11756
rect 28540 11704 28592 11756
rect 29276 11747 29328 11756
rect 29276 11713 29285 11747
rect 29285 11713 29319 11747
rect 29319 11713 29328 11747
rect 29276 11704 29328 11713
rect 30748 11747 30800 11756
rect 30748 11713 30757 11747
rect 30757 11713 30791 11747
rect 30791 11713 30800 11747
rect 30748 11704 30800 11713
rect 25872 11679 25924 11688
rect 25872 11645 25881 11679
rect 25881 11645 25915 11679
rect 25915 11645 25924 11679
rect 25872 11636 25924 11645
rect 26424 11636 26476 11688
rect 27160 11636 27212 11688
rect 26240 11568 26292 11620
rect 26516 11568 26568 11620
rect 27528 11636 27580 11688
rect 28724 11679 28776 11688
rect 28724 11645 28733 11679
rect 28733 11645 28767 11679
rect 28767 11645 28776 11679
rect 28724 11636 28776 11645
rect 30564 11636 30616 11688
rect 32496 11747 32548 11756
rect 24584 11543 24636 11552
rect 24584 11509 24593 11543
rect 24593 11509 24627 11543
rect 24627 11509 24636 11543
rect 24584 11500 24636 11509
rect 27252 11500 27304 11552
rect 31116 11568 31168 11620
rect 31300 11568 31352 11620
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 33048 11747 33100 11756
rect 33048 11713 33057 11747
rect 33057 11713 33091 11747
rect 33091 11713 33100 11747
rect 33048 11704 33100 11713
rect 33508 11636 33560 11688
rect 33968 11704 34020 11756
rect 34336 11772 34388 11824
rect 34244 11704 34296 11756
rect 35256 11772 35308 11824
rect 35624 11747 35676 11756
rect 35624 11713 35633 11747
rect 35633 11713 35667 11747
rect 35667 11713 35676 11747
rect 35624 11704 35676 11713
rect 36084 11747 36136 11756
rect 36084 11713 36093 11747
rect 36093 11713 36127 11747
rect 36127 11713 36136 11747
rect 36084 11704 36136 11713
rect 36636 11704 36688 11756
rect 36728 11747 36780 11756
rect 36728 11713 36737 11747
rect 36737 11713 36771 11747
rect 36771 11713 36780 11747
rect 36728 11704 36780 11713
rect 37188 11704 37240 11756
rect 37556 11840 37608 11892
rect 39028 11815 39080 11824
rect 39028 11781 39037 11815
rect 39037 11781 39071 11815
rect 39071 11781 39080 11815
rect 39028 11772 39080 11781
rect 39120 11772 39172 11824
rect 40224 11840 40276 11892
rect 40500 11840 40552 11892
rect 43260 11840 43312 11892
rect 44272 11883 44324 11892
rect 44272 11849 44281 11883
rect 44281 11849 44315 11883
rect 44315 11849 44324 11883
rect 44272 11840 44324 11849
rect 45560 11840 45612 11892
rect 37924 11747 37976 11756
rect 37924 11713 37933 11747
rect 37933 11713 37967 11747
rect 37967 11713 37976 11747
rect 37924 11704 37976 11713
rect 38660 11704 38712 11756
rect 40132 11704 40184 11756
rect 40316 11772 40368 11824
rect 43628 11772 43680 11824
rect 42340 11704 42392 11756
rect 42984 11747 43036 11756
rect 42984 11713 42993 11747
rect 42993 11713 43027 11747
rect 43027 11713 43036 11747
rect 42984 11704 43036 11713
rect 43076 11704 43128 11756
rect 43444 11747 43496 11756
rect 43444 11713 43453 11747
rect 43453 11713 43487 11747
rect 43487 11713 43496 11747
rect 43444 11704 43496 11713
rect 44456 11747 44508 11756
rect 44456 11713 44462 11747
rect 44462 11713 44496 11747
rect 44496 11713 44508 11747
rect 44916 11747 44968 11756
rect 44456 11704 44508 11713
rect 44916 11713 44925 11747
rect 44925 11713 44959 11747
rect 44959 11713 44968 11747
rect 44916 11704 44968 11713
rect 45560 11747 45612 11756
rect 45560 11713 45569 11747
rect 45569 11713 45603 11747
rect 45603 11713 45612 11747
rect 45560 11704 45612 11713
rect 45928 11840 45980 11892
rect 46296 11840 46348 11892
rect 46848 11883 46900 11892
rect 46848 11849 46857 11883
rect 46857 11849 46891 11883
rect 46891 11849 46900 11883
rect 46848 11840 46900 11849
rect 47400 11840 47452 11892
rect 47216 11772 47268 11824
rect 47768 11772 47820 11824
rect 48320 11883 48372 11892
rect 48320 11849 48329 11883
rect 48329 11849 48363 11883
rect 48363 11849 48372 11883
rect 48320 11840 48372 11849
rect 48504 11840 48556 11892
rect 49148 11840 49200 11892
rect 50620 11883 50672 11892
rect 50620 11849 50629 11883
rect 50629 11849 50663 11883
rect 50663 11849 50672 11883
rect 50620 11840 50672 11849
rect 50804 11883 50856 11892
rect 50804 11849 50813 11883
rect 50813 11849 50847 11883
rect 50847 11849 50856 11883
rect 50804 11840 50856 11849
rect 52000 11840 52052 11892
rect 48964 11772 49016 11824
rect 46112 11704 46164 11756
rect 46204 11704 46256 11756
rect 48596 11747 48648 11756
rect 32496 11568 32548 11620
rect 37004 11636 37056 11688
rect 27528 11500 27580 11552
rect 29828 11543 29880 11552
rect 29828 11509 29837 11543
rect 29837 11509 29871 11543
rect 29871 11509 29880 11543
rect 29828 11500 29880 11509
rect 31668 11500 31720 11552
rect 33232 11500 33284 11552
rect 33968 11500 34020 11552
rect 35348 11500 35400 11552
rect 36084 11500 36136 11552
rect 36728 11543 36780 11552
rect 36728 11509 36737 11543
rect 36737 11509 36771 11543
rect 36771 11509 36780 11543
rect 36728 11500 36780 11509
rect 37740 11636 37792 11688
rect 38476 11636 38528 11688
rect 42800 11636 42852 11688
rect 43996 11636 44048 11688
rect 37556 11568 37608 11620
rect 38936 11568 38988 11620
rect 45100 11568 45152 11620
rect 45652 11611 45704 11620
rect 37924 11500 37976 11552
rect 39212 11543 39264 11552
rect 39212 11509 39221 11543
rect 39221 11509 39255 11543
rect 39255 11509 39264 11543
rect 39212 11500 39264 11509
rect 40408 11500 40460 11552
rect 43352 11543 43404 11552
rect 43352 11509 43361 11543
rect 43361 11509 43395 11543
rect 43395 11509 43404 11543
rect 45652 11577 45661 11611
rect 45661 11577 45695 11611
rect 45695 11577 45704 11611
rect 45652 11568 45704 11577
rect 43352 11500 43404 11509
rect 46756 11500 46808 11552
rect 48596 11713 48605 11747
rect 48605 11713 48639 11747
rect 48639 11713 48648 11747
rect 48596 11704 48648 11713
rect 48688 11704 48740 11756
rect 48780 11636 48832 11688
rect 49148 11636 49200 11688
rect 49516 11679 49568 11688
rect 49516 11645 49525 11679
rect 49525 11645 49559 11679
rect 49559 11645 49568 11679
rect 49516 11636 49568 11645
rect 51080 11772 51132 11824
rect 51632 11636 51684 11688
rect 51356 11568 51408 11620
rect 48504 11500 48556 11552
rect 48780 11500 48832 11552
rect 49424 11543 49476 11552
rect 49424 11509 49433 11543
rect 49433 11509 49467 11543
rect 49467 11509 49476 11543
rect 49424 11500 49476 11509
rect 51724 11500 51776 11552
rect 52552 11840 52604 11892
rect 54208 11840 54260 11892
rect 55680 11840 55732 11892
rect 55956 11883 56008 11892
rect 55956 11849 55965 11883
rect 55965 11849 55999 11883
rect 55999 11849 56008 11883
rect 55956 11840 56008 11849
rect 53196 11772 53248 11824
rect 54484 11772 54536 11824
rect 52368 11747 52420 11756
rect 52368 11713 52377 11747
rect 52377 11713 52411 11747
rect 52411 11713 52420 11747
rect 52368 11704 52420 11713
rect 53564 11704 53616 11756
rect 54116 11747 54168 11756
rect 54116 11713 54125 11747
rect 54125 11713 54159 11747
rect 54159 11713 54168 11747
rect 54116 11704 54168 11713
rect 54576 11704 54628 11756
rect 55036 11747 55088 11756
rect 55036 11713 55045 11747
rect 55045 11713 55079 11747
rect 55079 11713 55088 11747
rect 55036 11704 55088 11713
rect 55496 11772 55548 11824
rect 55772 11815 55824 11824
rect 55772 11781 55797 11815
rect 55797 11781 55824 11815
rect 55772 11772 55824 11781
rect 53380 11636 53432 11688
rect 54208 11636 54260 11688
rect 52092 11568 52144 11620
rect 53288 11568 53340 11620
rect 54852 11611 54904 11620
rect 54852 11577 54861 11611
rect 54861 11577 54895 11611
rect 54895 11577 54904 11611
rect 54852 11568 54904 11577
rect 52736 11500 52788 11552
rect 55680 11500 55732 11552
rect 57428 11500 57480 11552
rect 57888 11500 57940 11552
rect 58256 11500 58308 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 26056 11296 26108 11348
rect 27436 11339 27488 11348
rect 27436 11305 27445 11339
rect 27445 11305 27479 11339
rect 27479 11305 27488 11339
rect 27436 11296 27488 11305
rect 28264 11339 28316 11348
rect 28264 11305 28273 11339
rect 28273 11305 28307 11339
rect 28307 11305 28316 11339
rect 28264 11296 28316 11305
rect 28816 11296 28868 11348
rect 29000 11296 29052 11348
rect 25688 11228 25740 11280
rect 27344 11228 27396 11280
rect 28908 11228 28960 11280
rect 29460 11228 29512 11280
rect 30656 11296 30708 11348
rect 32312 11296 32364 11348
rect 32956 11339 33008 11348
rect 32956 11305 32965 11339
rect 32965 11305 32999 11339
rect 32999 11305 33008 11339
rect 32956 11296 33008 11305
rect 33784 11296 33836 11348
rect 33968 11296 34020 11348
rect 35624 11296 35676 11348
rect 35900 11296 35952 11348
rect 36360 11296 36412 11348
rect 37740 11339 37792 11348
rect 37740 11305 37749 11339
rect 37749 11305 37783 11339
rect 37783 11305 37792 11339
rect 37740 11296 37792 11305
rect 37924 11296 37976 11348
rect 38568 11296 38620 11348
rect 40776 11339 40828 11348
rect 40776 11305 40785 11339
rect 40785 11305 40819 11339
rect 40819 11305 40828 11339
rect 40776 11296 40828 11305
rect 42340 11339 42392 11348
rect 42340 11305 42349 11339
rect 42349 11305 42383 11339
rect 42383 11305 42392 11339
rect 42340 11296 42392 11305
rect 43352 11296 43404 11348
rect 43996 11339 44048 11348
rect 43996 11305 44005 11339
rect 44005 11305 44039 11339
rect 44039 11305 44048 11339
rect 43996 11296 44048 11305
rect 33508 11228 33560 11280
rect 27896 11160 27948 11212
rect 30288 11160 30340 11212
rect 31668 11160 31720 11212
rect 23848 11024 23900 11076
rect 25044 11092 25096 11144
rect 25964 11092 26016 11144
rect 28172 11092 28224 11144
rect 28356 11092 28408 11144
rect 26148 11024 26200 11076
rect 27620 11067 27672 11076
rect 27620 11033 27629 11067
rect 27629 11033 27663 11067
rect 27663 11033 27672 11067
rect 27620 11024 27672 11033
rect 28264 11024 28316 11076
rect 28908 11092 28960 11144
rect 29460 11024 29512 11076
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 30564 11092 30616 11144
rect 30932 11135 30984 11144
rect 30932 11101 30941 11135
rect 30941 11101 30975 11135
rect 30975 11101 30984 11135
rect 30932 11092 30984 11101
rect 31208 11092 31260 11144
rect 32036 11135 32088 11144
rect 32036 11101 32045 11135
rect 32045 11101 32079 11135
rect 32079 11101 32088 11135
rect 32036 11092 32088 11101
rect 33048 11160 33100 11212
rect 34888 11228 34940 11280
rect 35808 11228 35860 11280
rect 36544 11271 36596 11280
rect 36544 11237 36553 11271
rect 36553 11237 36587 11271
rect 36587 11237 36596 11271
rect 36544 11228 36596 11237
rect 37280 11228 37332 11280
rect 38108 11228 38160 11280
rect 39396 11228 39448 11280
rect 43720 11228 43772 11280
rect 46940 11296 46992 11348
rect 47768 11296 47820 11348
rect 48688 11296 48740 11348
rect 49056 11296 49108 11348
rect 45100 11228 45152 11280
rect 45928 11228 45980 11280
rect 47216 11228 47268 11280
rect 50712 11228 50764 11280
rect 35624 11160 35676 11212
rect 29828 11024 29880 11076
rect 25688 10956 25740 11008
rect 26884 10999 26936 11008
rect 26884 10965 26893 10999
rect 26893 10965 26927 10999
rect 26927 10965 26936 10999
rect 26884 10956 26936 10965
rect 27252 10956 27304 11008
rect 31208 10956 31260 11008
rect 31392 11024 31444 11076
rect 34428 11092 34480 11144
rect 35532 11135 35584 11144
rect 35532 11101 35541 11135
rect 35541 11101 35575 11135
rect 35575 11101 35584 11135
rect 36820 11135 36872 11144
rect 35532 11092 35584 11101
rect 36820 11101 36829 11135
rect 36829 11101 36863 11135
rect 36863 11101 36872 11135
rect 36820 11092 36872 11101
rect 37188 11092 37240 11144
rect 37556 11135 37608 11144
rect 37556 11101 37565 11135
rect 37565 11101 37599 11135
rect 37599 11101 37608 11135
rect 37556 11092 37608 11101
rect 38660 11160 38712 11212
rect 42708 11160 42760 11212
rect 43168 11160 43220 11212
rect 39028 11092 39080 11144
rect 40408 11135 40460 11144
rect 40408 11101 40417 11135
rect 40417 11101 40451 11135
rect 40451 11101 40460 11135
rect 40408 11092 40460 11101
rect 42616 11092 42668 11144
rect 32772 11067 32824 11076
rect 32772 11033 32781 11067
rect 32781 11033 32815 11067
rect 32815 11033 32824 11067
rect 32772 11024 32824 11033
rect 32956 11067 33008 11076
rect 32956 11033 32965 11067
rect 32965 11033 32999 11067
rect 32999 11033 33008 11067
rect 32956 11024 33008 11033
rect 34244 11024 34296 11076
rect 36912 11024 36964 11076
rect 31668 10956 31720 11008
rect 35440 10956 35492 11008
rect 37372 10999 37424 11008
rect 37372 10965 37381 10999
rect 37381 10965 37415 10999
rect 37415 10965 37424 10999
rect 40224 11024 40276 11076
rect 41788 10999 41840 11008
rect 37372 10956 37424 10965
rect 41788 10965 41797 10999
rect 41797 10965 41831 10999
rect 41831 10965 41840 10999
rect 41788 10956 41840 10965
rect 44824 11092 44876 11144
rect 45560 11160 45612 11212
rect 47492 11203 47544 11212
rect 47492 11169 47501 11203
rect 47501 11169 47535 11203
rect 47535 11169 47544 11203
rect 47492 11160 47544 11169
rect 47308 11135 47360 11144
rect 47308 11101 47317 11135
rect 47317 11101 47351 11135
rect 47351 11101 47360 11135
rect 47308 11092 47360 11101
rect 47584 11135 47636 11144
rect 47584 11101 47593 11135
rect 47593 11101 47627 11135
rect 47627 11101 47636 11135
rect 47584 11092 47636 11101
rect 43168 11024 43220 11076
rect 44548 11067 44600 11076
rect 44548 11033 44557 11067
rect 44557 11033 44591 11067
rect 44591 11033 44600 11067
rect 44548 11024 44600 11033
rect 45744 11024 45796 11076
rect 47400 11024 47452 11076
rect 47768 11092 47820 11144
rect 48320 11135 48372 11144
rect 48320 11101 48329 11135
rect 48329 11101 48363 11135
rect 48363 11101 48372 11135
rect 48504 11135 48556 11144
rect 48320 11092 48372 11101
rect 48504 11101 48513 11135
rect 48513 11101 48547 11135
rect 48547 11101 48556 11135
rect 48504 11092 48556 11101
rect 48780 11092 48832 11144
rect 49976 11092 50028 11144
rect 50160 11092 50212 11144
rect 50528 11135 50580 11144
rect 50528 11101 50537 11135
rect 50537 11101 50571 11135
rect 50571 11101 50580 11135
rect 50528 11092 50580 11101
rect 50896 11296 50948 11348
rect 52184 11296 52236 11348
rect 54208 11296 54260 11348
rect 54300 11296 54352 11348
rect 55772 11296 55824 11348
rect 58072 11339 58124 11348
rect 51080 11228 51132 11280
rect 53748 11160 53800 11212
rect 54484 11160 54536 11212
rect 49700 11024 49752 11076
rect 50068 11024 50120 11076
rect 51080 11092 51132 11144
rect 51540 11092 51592 11144
rect 52000 11135 52052 11144
rect 52000 11101 52009 11135
rect 52009 11101 52043 11135
rect 52043 11101 52052 11135
rect 52000 11092 52052 11101
rect 51632 11024 51684 11076
rect 52092 11024 52144 11076
rect 53012 11092 53064 11144
rect 53104 11092 53156 11144
rect 53288 11024 53340 11076
rect 54116 11135 54168 11144
rect 54116 11101 54125 11135
rect 54125 11101 54159 11135
rect 54159 11101 54168 11135
rect 54116 11092 54168 11101
rect 55036 11092 55088 11144
rect 54392 11024 54444 11076
rect 54852 11067 54904 11076
rect 54852 11033 54861 11067
rect 54861 11033 54895 11067
rect 54895 11033 54904 11067
rect 54852 11024 54904 11033
rect 43996 10956 44048 11008
rect 44088 10956 44140 11008
rect 45928 10956 45980 11008
rect 48044 10956 48096 11008
rect 48228 10956 48280 11008
rect 50528 10956 50580 11008
rect 50712 10956 50764 11008
rect 50896 10956 50948 11008
rect 52552 10956 52604 11008
rect 53104 10956 53156 11008
rect 53564 10956 53616 11008
rect 55312 11024 55364 11076
rect 55680 11067 55732 11076
rect 55680 11033 55689 11067
rect 55689 11033 55723 11067
rect 55723 11033 55732 11067
rect 55680 11024 55732 11033
rect 58072 11305 58081 11339
rect 58081 11305 58115 11339
rect 58115 11305 58124 11339
rect 58072 11296 58124 11305
rect 55772 10956 55824 11008
rect 56508 10956 56560 11008
rect 56692 10956 56744 11008
rect 57520 10999 57572 11008
rect 57520 10965 57529 10999
rect 57529 10965 57563 10999
rect 57563 10965 57572 10999
rect 57520 10956 57572 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 24492 10752 24544 10804
rect 25228 10684 25280 10736
rect 24768 10616 24820 10668
rect 26424 10684 26476 10736
rect 27436 10684 27488 10736
rect 27344 10659 27396 10668
rect 27344 10625 27353 10659
rect 27353 10625 27387 10659
rect 27387 10625 27396 10659
rect 27344 10616 27396 10625
rect 27620 10659 27672 10668
rect 27620 10625 27629 10659
rect 27629 10625 27663 10659
rect 27663 10625 27672 10659
rect 27620 10616 27672 10625
rect 28632 10727 28684 10736
rect 28632 10693 28641 10727
rect 28641 10693 28675 10727
rect 28675 10693 28684 10727
rect 28632 10684 28684 10693
rect 29460 10752 29512 10804
rect 29920 10752 29972 10804
rect 30288 10795 30340 10804
rect 30288 10761 30297 10795
rect 30297 10761 30331 10795
rect 30331 10761 30340 10795
rect 30288 10752 30340 10761
rect 30380 10752 30432 10804
rect 30748 10752 30800 10804
rect 30932 10752 30984 10804
rect 31300 10752 31352 10804
rect 32036 10752 32088 10804
rect 33692 10752 33744 10804
rect 34612 10752 34664 10804
rect 35348 10752 35400 10804
rect 29184 10616 29236 10668
rect 24676 10591 24728 10600
rect 24676 10557 24685 10591
rect 24685 10557 24719 10591
rect 24719 10557 24728 10591
rect 24676 10548 24728 10557
rect 26976 10548 27028 10600
rect 27344 10480 27396 10532
rect 28816 10591 28868 10600
rect 28816 10557 28825 10591
rect 28825 10557 28859 10591
rect 28859 10557 28868 10591
rect 28816 10548 28868 10557
rect 24860 10455 24912 10464
rect 24860 10421 24869 10455
rect 24869 10421 24903 10455
rect 24903 10421 24912 10455
rect 24860 10412 24912 10421
rect 25228 10412 25280 10464
rect 26516 10412 26568 10464
rect 26792 10412 26844 10464
rect 27252 10412 27304 10464
rect 29276 10480 29328 10532
rect 29920 10659 29972 10668
rect 29920 10625 29929 10659
rect 29929 10625 29963 10659
rect 29963 10625 29972 10659
rect 30104 10659 30156 10668
rect 29920 10616 29972 10625
rect 30104 10625 30127 10659
rect 30127 10625 30156 10659
rect 30104 10616 30156 10625
rect 32772 10684 32824 10736
rect 33048 10684 33100 10736
rect 31760 10616 31812 10668
rect 33876 10616 33928 10668
rect 34612 10616 34664 10668
rect 38384 10752 38436 10804
rect 40224 10752 40276 10804
rect 36360 10684 36412 10736
rect 37648 10684 37700 10736
rect 30196 10548 30248 10600
rect 32220 10480 32272 10532
rect 32588 10480 32640 10532
rect 32772 10591 32824 10600
rect 32772 10557 32781 10591
rect 32781 10557 32815 10591
rect 32815 10557 32824 10591
rect 32772 10548 32824 10557
rect 34244 10591 34296 10600
rect 34244 10557 34253 10591
rect 34253 10557 34287 10591
rect 34287 10557 34296 10591
rect 34244 10548 34296 10557
rect 34336 10591 34388 10600
rect 34336 10557 34345 10591
rect 34345 10557 34379 10591
rect 34379 10557 34388 10591
rect 35256 10591 35308 10600
rect 34336 10548 34388 10557
rect 35256 10557 35265 10591
rect 35265 10557 35299 10591
rect 35299 10557 35308 10591
rect 35256 10548 35308 10557
rect 36452 10616 36504 10668
rect 35900 10548 35952 10600
rect 37280 10616 37332 10668
rect 37832 10684 37884 10736
rect 38568 10659 38620 10668
rect 38568 10625 38577 10659
rect 38577 10625 38611 10659
rect 38611 10625 38620 10659
rect 38568 10616 38620 10625
rect 38936 10616 38988 10668
rect 39396 10659 39448 10668
rect 39396 10625 39405 10659
rect 39405 10625 39439 10659
rect 39439 10625 39448 10659
rect 39396 10616 39448 10625
rect 40684 10659 40736 10668
rect 40684 10625 40693 10659
rect 40693 10625 40727 10659
rect 40727 10625 40736 10659
rect 41788 10684 41840 10736
rect 42340 10684 42392 10736
rect 43444 10684 43496 10736
rect 44088 10684 44140 10736
rect 40684 10616 40736 10625
rect 42432 10616 42484 10668
rect 44272 10659 44324 10668
rect 44272 10625 44281 10659
rect 44281 10625 44315 10659
rect 44315 10625 44324 10659
rect 44272 10616 44324 10625
rect 45560 10684 45612 10736
rect 46848 10752 46900 10804
rect 46112 10659 46164 10668
rect 46112 10625 46121 10659
rect 46121 10625 46155 10659
rect 46155 10625 46164 10659
rect 46112 10616 46164 10625
rect 46296 10616 46348 10668
rect 46664 10616 46716 10668
rect 38292 10548 38344 10600
rect 38476 10591 38528 10600
rect 38476 10557 38485 10591
rect 38485 10557 38519 10591
rect 38519 10557 38528 10591
rect 38476 10548 38528 10557
rect 39304 10548 39356 10600
rect 39764 10548 39816 10600
rect 45652 10548 45704 10600
rect 46572 10548 46624 10600
rect 48044 10727 48096 10736
rect 48044 10693 48053 10727
rect 48053 10693 48087 10727
rect 48087 10693 48096 10727
rect 48044 10684 48096 10693
rect 51080 10752 51132 10804
rect 47768 10659 47820 10668
rect 47768 10625 47777 10659
rect 47777 10625 47811 10659
rect 47811 10625 47820 10659
rect 47768 10616 47820 10625
rect 48872 10659 48924 10668
rect 48872 10625 48881 10659
rect 48881 10625 48915 10659
rect 48915 10625 48924 10659
rect 48872 10616 48924 10625
rect 49700 10591 49752 10600
rect 28080 10412 28132 10464
rect 28540 10412 28592 10464
rect 30932 10412 30984 10464
rect 31208 10455 31260 10464
rect 31208 10421 31226 10455
rect 31226 10421 31260 10455
rect 46480 10523 46532 10532
rect 46480 10489 46489 10523
rect 46489 10489 46523 10523
rect 46523 10489 46532 10523
rect 46480 10480 46532 10489
rect 46664 10480 46716 10532
rect 49700 10557 49709 10591
rect 49709 10557 49743 10591
rect 49743 10557 49752 10591
rect 49700 10548 49752 10557
rect 47032 10480 47084 10532
rect 49516 10480 49568 10532
rect 50160 10616 50212 10668
rect 51724 10684 51776 10736
rect 52000 10752 52052 10804
rect 54024 10795 54076 10804
rect 54024 10761 54033 10795
rect 54033 10761 54067 10795
rect 54067 10761 54076 10795
rect 54024 10752 54076 10761
rect 54208 10752 54260 10804
rect 53012 10727 53064 10736
rect 51632 10659 51684 10668
rect 51632 10625 51641 10659
rect 51641 10625 51675 10659
rect 51675 10625 51684 10659
rect 51632 10616 51684 10625
rect 52092 10659 52144 10668
rect 52092 10625 52101 10659
rect 52101 10625 52135 10659
rect 52135 10625 52144 10659
rect 52092 10616 52144 10625
rect 52184 10616 52236 10668
rect 50528 10591 50580 10600
rect 50528 10557 50537 10591
rect 50537 10557 50571 10591
rect 50571 10557 50580 10591
rect 50528 10548 50580 10557
rect 51356 10548 51408 10600
rect 52460 10548 52512 10600
rect 53012 10693 53021 10727
rect 53021 10693 53055 10727
rect 53055 10693 53064 10727
rect 55128 10752 55180 10804
rect 58256 10752 58308 10804
rect 53012 10684 53064 10693
rect 55496 10684 55548 10736
rect 56324 10684 56376 10736
rect 52920 10659 52972 10668
rect 52920 10625 52929 10659
rect 52929 10625 52963 10659
rect 52963 10625 52972 10659
rect 52920 10616 52972 10625
rect 53288 10616 53340 10668
rect 54208 10659 54260 10668
rect 54208 10625 54217 10659
rect 54217 10625 54251 10659
rect 54251 10625 54260 10659
rect 54208 10616 54260 10625
rect 54300 10659 54352 10668
rect 54300 10625 54309 10659
rect 54309 10625 54343 10659
rect 54343 10625 54352 10659
rect 54576 10659 54628 10668
rect 54300 10616 54352 10625
rect 54576 10625 54585 10659
rect 54585 10625 54619 10659
rect 54619 10625 54628 10659
rect 54576 10616 54628 10625
rect 56140 10616 56192 10668
rect 54484 10591 54536 10600
rect 54484 10557 54493 10591
rect 54493 10557 54527 10591
rect 54527 10557 54536 10591
rect 54484 10548 54536 10557
rect 31208 10412 31260 10421
rect 35532 10412 35584 10464
rect 36728 10455 36780 10464
rect 36728 10421 36737 10455
rect 36737 10421 36771 10455
rect 36771 10421 36780 10455
rect 36728 10412 36780 10421
rect 43076 10412 43128 10464
rect 43720 10412 43772 10464
rect 44088 10455 44140 10464
rect 44088 10421 44097 10455
rect 44097 10421 44131 10455
rect 44131 10421 44140 10455
rect 44088 10412 44140 10421
rect 45376 10455 45428 10464
rect 45376 10421 45385 10455
rect 45385 10421 45419 10455
rect 45419 10421 45428 10455
rect 45376 10412 45428 10421
rect 45836 10412 45888 10464
rect 46940 10412 46992 10464
rect 49424 10412 49476 10464
rect 49792 10455 49844 10464
rect 49792 10421 49801 10455
rect 49801 10421 49835 10455
rect 49835 10421 49844 10455
rect 49792 10412 49844 10421
rect 51356 10412 51408 10464
rect 52644 10412 52696 10464
rect 55312 10412 55364 10464
rect 56784 10455 56836 10464
rect 56784 10421 56793 10455
rect 56793 10421 56827 10455
rect 56827 10421 56836 10455
rect 56784 10412 56836 10421
rect 57980 10412 58032 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 24676 10208 24728 10260
rect 26332 10208 26384 10260
rect 26792 10251 26844 10260
rect 26792 10217 26801 10251
rect 26801 10217 26835 10251
rect 26835 10217 26844 10251
rect 26792 10208 26844 10217
rect 27712 10208 27764 10260
rect 27988 10208 28040 10260
rect 28448 10251 28500 10260
rect 28448 10217 28457 10251
rect 28457 10217 28491 10251
rect 28491 10217 28500 10251
rect 28448 10208 28500 10217
rect 28632 10208 28684 10260
rect 28908 10208 28960 10260
rect 29184 10251 29236 10260
rect 29184 10217 29193 10251
rect 29193 10217 29227 10251
rect 29227 10217 29236 10251
rect 29184 10208 29236 10217
rect 29828 10208 29880 10260
rect 30196 10208 30248 10260
rect 30564 10251 30616 10260
rect 30564 10217 30573 10251
rect 30573 10217 30607 10251
rect 30607 10217 30616 10251
rect 30564 10208 30616 10217
rect 31760 10208 31812 10260
rect 33140 10208 33192 10260
rect 33784 10208 33836 10260
rect 36452 10208 36504 10260
rect 37556 10208 37608 10260
rect 38660 10208 38712 10260
rect 38752 10208 38804 10260
rect 28540 10140 28592 10192
rect 23848 10047 23900 10056
rect 23848 10013 23857 10047
rect 23857 10013 23891 10047
rect 23891 10013 23900 10047
rect 23848 10004 23900 10013
rect 25228 10072 25280 10124
rect 27160 10072 27212 10124
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 24584 9979 24636 9988
rect 24584 9945 24593 9979
rect 24593 9945 24627 9979
rect 24627 9945 24636 9979
rect 24584 9936 24636 9945
rect 24768 9979 24820 9988
rect 24768 9945 24777 9979
rect 24777 9945 24811 9979
rect 24811 9945 24820 9979
rect 24768 9936 24820 9945
rect 25964 10004 26016 10056
rect 26608 10004 26660 10056
rect 26884 10047 26936 10056
rect 26884 10013 26893 10047
rect 26893 10013 26927 10047
rect 26927 10013 26936 10047
rect 26884 10004 26936 10013
rect 27344 10004 27396 10056
rect 26332 9936 26384 9988
rect 28080 10047 28132 10056
rect 28080 10013 28089 10047
rect 28089 10013 28123 10047
rect 28123 10013 28132 10047
rect 28080 10004 28132 10013
rect 28816 10004 28868 10056
rect 29092 10004 29144 10056
rect 29828 10004 29880 10056
rect 30104 10004 30156 10056
rect 30564 10047 30616 10056
rect 30564 10013 30573 10047
rect 30573 10013 30607 10047
rect 30607 10013 30616 10047
rect 30564 10004 30616 10013
rect 31300 10004 31352 10056
rect 32772 10072 32824 10124
rect 33876 10115 33928 10124
rect 31668 10047 31720 10056
rect 31208 9936 31260 9988
rect 31668 10013 31677 10047
rect 31677 10013 31711 10047
rect 31711 10013 31720 10047
rect 31668 10004 31720 10013
rect 32220 10004 32272 10056
rect 33876 10081 33885 10115
rect 33885 10081 33919 10115
rect 33919 10081 33928 10115
rect 33876 10072 33928 10081
rect 33968 10072 34020 10124
rect 31944 9936 31996 9988
rect 25688 9911 25740 9920
rect 25688 9877 25697 9911
rect 25697 9877 25731 9911
rect 25731 9877 25740 9911
rect 25688 9868 25740 9877
rect 28356 9868 28408 9920
rect 29552 9868 29604 9920
rect 29920 9868 29972 9920
rect 30104 9868 30156 9920
rect 31300 9868 31352 9920
rect 31668 9868 31720 9920
rect 32772 9868 32824 9920
rect 33232 10047 33284 10056
rect 33232 10013 33253 10047
rect 33253 10013 33284 10047
rect 33232 10004 33284 10013
rect 34060 10047 34112 10056
rect 33508 9936 33560 9988
rect 33692 9979 33744 9988
rect 33692 9945 33701 9979
rect 33701 9945 33735 9979
rect 33735 9945 33744 9979
rect 33692 9936 33744 9945
rect 34060 10013 34069 10047
rect 34069 10013 34103 10047
rect 34103 10013 34112 10047
rect 34060 10004 34112 10013
rect 35992 10140 36044 10192
rect 34336 10072 34388 10124
rect 36544 10115 36596 10124
rect 35808 10047 35860 10056
rect 35808 10013 35817 10047
rect 35817 10013 35851 10047
rect 35851 10013 35860 10047
rect 35808 10004 35860 10013
rect 36544 10081 36553 10115
rect 36553 10081 36587 10115
rect 36587 10081 36596 10115
rect 36544 10072 36596 10081
rect 41236 10072 41288 10124
rect 36912 10047 36964 10056
rect 36176 9936 36228 9988
rect 34336 9868 34388 9920
rect 34612 9868 34664 9920
rect 34796 9868 34848 9920
rect 35808 9868 35860 9920
rect 36912 10013 36921 10047
rect 36921 10013 36955 10047
rect 36955 10013 36964 10047
rect 36912 10004 36964 10013
rect 38844 10004 38896 10056
rect 39120 10047 39172 10056
rect 39120 10013 39129 10047
rect 39129 10013 39163 10047
rect 39163 10013 39172 10047
rect 39120 10004 39172 10013
rect 39212 10047 39264 10056
rect 39212 10013 39221 10047
rect 39221 10013 39255 10047
rect 39255 10013 39264 10047
rect 39212 10004 39264 10013
rect 40224 10047 40276 10056
rect 40224 10013 40233 10047
rect 40233 10013 40267 10047
rect 40267 10013 40276 10047
rect 40224 10004 40276 10013
rect 41328 10047 41380 10056
rect 41328 10013 41337 10047
rect 41337 10013 41371 10047
rect 41371 10013 41380 10047
rect 41328 10004 41380 10013
rect 45652 10208 45704 10260
rect 45928 10251 45980 10260
rect 45928 10217 45937 10251
rect 45937 10217 45971 10251
rect 45971 10217 45980 10251
rect 45928 10208 45980 10217
rect 46112 10208 46164 10260
rect 47676 10251 47728 10260
rect 47676 10217 47685 10251
rect 47685 10217 47719 10251
rect 47719 10217 47728 10251
rect 47676 10208 47728 10217
rect 49240 10208 49292 10260
rect 49424 10208 49476 10260
rect 50436 10208 50488 10260
rect 51632 10208 51684 10260
rect 52184 10208 52236 10260
rect 52644 10208 52696 10260
rect 53104 10208 53156 10260
rect 53748 10208 53800 10260
rect 54116 10208 54168 10260
rect 45376 10183 45428 10192
rect 45376 10149 45385 10183
rect 45385 10149 45419 10183
rect 45419 10149 45428 10183
rect 45376 10140 45428 10149
rect 48872 10140 48924 10192
rect 44088 10004 44140 10056
rect 44364 10004 44416 10056
rect 36544 9936 36596 9988
rect 37004 9936 37056 9988
rect 38108 9979 38160 9988
rect 38108 9945 38117 9979
rect 38117 9945 38151 9979
rect 38151 9945 38160 9979
rect 38108 9936 38160 9945
rect 38292 9979 38344 9988
rect 38292 9945 38317 9979
rect 38317 9945 38344 9979
rect 40408 9979 40460 9988
rect 38292 9936 38344 9945
rect 40408 9945 40417 9979
rect 40417 9945 40451 9979
rect 40451 9945 40460 9979
rect 40408 9936 40460 9945
rect 43168 9936 43220 9988
rect 43352 9979 43404 9988
rect 43352 9945 43361 9979
rect 43361 9945 43395 9979
rect 43395 9945 43404 9979
rect 43352 9936 43404 9945
rect 43996 9979 44048 9988
rect 43996 9945 44023 9979
rect 44023 9945 44048 9979
rect 43996 9936 44048 9945
rect 44548 9936 44600 9988
rect 46756 10072 46808 10124
rect 45744 10047 45796 10056
rect 45744 10013 45756 10047
rect 45756 10013 45790 10047
rect 45790 10013 45796 10047
rect 45744 10004 45796 10013
rect 46848 10047 46900 10056
rect 46848 10013 46857 10047
rect 46857 10013 46891 10047
rect 46891 10013 46900 10047
rect 46848 10004 46900 10013
rect 48688 10072 48740 10124
rect 50160 10140 50212 10192
rect 50896 10140 50948 10192
rect 51448 10183 51500 10192
rect 51448 10149 51457 10183
rect 51457 10149 51491 10183
rect 51491 10149 51500 10183
rect 51448 10140 51500 10149
rect 51540 10183 51592 10192
rect 51540 10149 51549 10183
rect 51549 10149 51583 10183
rect 51583 10149 51592 10183
rect 51540 10140 51592 10149
rect 51724 10140 51776 10192
rect 52000 10140 52052 10192
rect 48136 10047 48188 10056
rect 45928 9936 45980 9988
rect 46204 9936 46256 9988
rect 46756 9936 46808 9988
rect 43444 9868 43496 9920
rect 45744 9911 45796 9920
rect 45744 9877 45753 9911
rect 45753 9877 45787 9911
rect 45787 9877 45796 9911
rect 45744 9868 45796 9877
rect 48136 10013 48145 10047
rect 48145 10013 48179 10047
rect 48179 10013 48188 10047
rect 48136 10004 48188 10013
rect 49056 10004 49108 10056
rect 49424 10047 49476 10056
rect 49424 10013 49433 10047
rect 49433 10013 49467 10047
rect 49467 10013 49476 10047
rect 49424 10004 49476 10013
rect 53012 10072 53064 10124
rect 53288 10140 53340 10192
rect 56692 10208 56744 10260
rect 55680 10140 55732 10192
rect 50436 10004 50488 10056
rect 50804 10047 50856 10056
rect 50804 10013 50813 10047
rect 50813 10013 50847 10047
rect 50847 10013 50856 10047
rect 50804 10004 50856 10013
rect 51356 10047 51408 10056
rect 51356 10013 51365 10047
rect 51365 10013 51399 10047
rect 51399 10013 51408 10047
rect 51356 10004 51408 10013
rect 51632 10047 51684 10056
rect 51632 10013 51641 10047
rect 51641 10013 51675 10047
rect 51675 10013 51684 10047
rect 51632 10004 51684 10013
rect 53104 10047 53156 10056
rect 53104 10013 53113 10047
rect 53113 10013 53147 10047
rect 53147 10013 53156 10047
rect 53104 10004 53156 10013
rect 56784 10072 56836 10124
rect 53748 10047 53800 10056
rect 53748 10013 53757 10047
rect 53757 10013 53791 10047
rect 53791 10013 53800 10047
rect 53748 10004 53800 10013
rect 56140 10047 56192 10056
rect 49792 9979 49844 9988
rect 49792 9945 49801 9979
rect 49801 9945 49835 9979
rect 49835 9945 49844 9979
rect 49792 9936 49844 9945
rect 53840 9936 53892 9988
rect 50712 9868 50764 9920
rect 53104 9868 53156 9920
rect 53472 9868 53524 9920
rect 53748 9868 53800 9920
rect 56140 10013 56149 10047
rect 56149 10013 56183 10047
rect 56183 10013 56192 10047
rect 56140 10004 56192 10013
rect 56416 10047 56468 10056
rect 56416 10013 56425 10047
rect 56425 10013 56459 10047
rect 56459 10013 56468 10047
rect 56416 10004 56468 10013
rect 57244 10004 57296 10056
rect 57980 10004 58032 10056
rect 55312 9868 55364 9920
rect 57428 9936 57480 9988
rect 56968 9868 57020 9920
rect 57152 9868 57204 9920
rect 57612 9911 57664 9920
rect 57612 9877 57621 9911
rect 57621 9877 57655 9911
rect 57655 9877 57664 9911
rect 57612 9868 57664 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 26884 9664 26936 9716
rect 28816 9664 28868 9716
rect 24124 9596 24176 9648
rect 25780 9596 25832 9648
rect 26792 9596 26844 9648
rect 27252 9596 27304 9648
rect 27804 9596 27856 9648
rect 28356 9596 28408 9648
rect 28540 9596 28592 9648
rect 25964 9528 26016 9580
rect 27896 9528 27948 9580
rect 28264 9528 28316 9580
rect 28632 9571 28684 9580
rect 28632 9537 28641 9571
rect 28641 9537 28675 9571
rect 28675 9537 28684 9571
rect 28632 9528 28684 9537
rect 24584 9460 24636 9512
rect 26608 9460 26660 9512
rect 27620 9460 27672 9512
rect 28816 9460 28868 9512
rect 29552 9528 29604 9580
rect 29828 9571 29880 9580
rect 29828 9537 29837 9571
rect 29837 9537 29871 9571
rect 29871 9537 29880 9571
rect 29828 9528 29880 9537
rect 30104 9571 30156 9580
rect 30104 9537 30113 9571
rect 30113 9537 30147 9571
rect 30147 9537 30156 9571
rect 30104 9528 30156 9537
rect 31116 9596 31168 9648
rect 30932 9571 30984 9580
rect 30932 9537 30941 9571
rect 30941 9537 30975 9571
rect 30975 9537 30984 9571
rect 30932 9528 30984 9537
rect 31208 9571 31260 9580
rect 30012 9460 30064 9512
rect 30564 9460 30616 9512
rect 31208 9537 31217 9571
rect 31217 9537 31251 9571
rect 31251 9537 31260 9571
rect 31208 9528 31260 9537
rect 33876 9664 33928 9716
rect 31576 9596 31628 9648
rect 32404 9596 32456 9648
rect 32680 9596 32732 9648
rect 32956 9571 33008 9614
rect 32956 9562 32982 9571
rect 32982 9562 33008 9571
rect 34060 9596 34112 9648
rect 33048 9571 33100 9580
rect 33048 9537 33057 9571
rect 33057 9537 33091 9571
rect 33091 9537 33100 9571
rect 33324 9571 33376 9580
rect 33048 9528 33100 9537
rect 33324 9537 33333 9571
rect 33333 9537 33367 9571
rect 33367 9537 33376 9571
rect 33324 9528 33376 9537
rect 33876 9528 33928 9580
rect 32036 9460 32088 9512
rect 29368 9392 29420 9444
rect 29644 9392 29696 9444
rect 24952 9367 25004 9376
rect 24952 9333 24961 9367
rect 24961 9333 24995 9367
rect 24995 9333 25004 9367
rect 24952 9324 25004 9333
rect 26424 9324 26476 9376
rect 27252 9324 27304 9376
rect 27712 9324 27764 9376
rect 28356 9324 28408 9376
rect 30104 9392 30156 9444
rect 30656 9392 30708 9444
rect 31116 9392 31168 9444
rect 33140 9392 33192 9444
rect 33508 9392 33560 9444
rect 31300 9324 31352 9376
rect 34060 9324 34112 9376
rect 36176 9639 36228 9648
rect 36176 9605 36201 9639
rect 36201 9605 36228 9639
rect 36912 9664 36964 9716
rect 39764 9707 39816 9716
rect 36176 9596 36228 9605
rect 36544 9528 36596 9580
rect 37280 9528 37332 9580
rect 39764 9673 39773 9707
rect 39773 9673 39807 9707
rect 39807 9673 39816 9707
rect 39764 9664 39816 9673
rect 44272 9664 44324 9716
rect 45468 9664 45520 9716
rect 46480 9664 46532 9716
rect 48596 9664 48648 9716
rect 49332 9664 49384 9716
rect 52092 9664 52144 9716
rect 56140 9664 56192 9716
rect 56416 9664 56468 9716
rect 39396 9596 39448 9648
rect 44364 9639 44416 9648
rect 44364 9605 44373 9639
rect 44373 9605 44407 9639
rect 44407 9605 44416 9639
rect 44364 9596 44416 9605
rect 45928 9596 45980 9648
rect 47124 9596 47176 9648
rect 48688 9639 48740 9648
rect 48688 9605 48697 9639
rect 48697 9605 48731 9639
rect 48731 9605 48740 9639
rect 48688 9596 48740 9605
rect 35440 9460 35492 9512
rect 37004 9460 37056 9512
rect 38108 9528 38160 9580
rect 39580 9571 39632 9580
rect 39580 9537 39589 9571
rect 39589 9537 39623 9571
rect 39623 9537 39632 9571
rect 39580 9528 39632 9537
rect 40224 9528 40276 9580
rect 41236 9528 41288 9580
rect 38752 9460 38804 9512
rect 34428 9392 34480 9444
rect 38108 9392 38160 9444
rect 38200 9392 38252 9444
rect 40960 9392 41012 9444
rect 43996 9528 44048 9580
rect 44732 9528 44784 9580
rect 45284 9528 45336 9580
rect 45836 9571 45888 9580
rect 45836 9537 45845 9571
rect 45845 9537 45879 9571
rect 45879 9537 45888 9571
rect 45836 9528 45888 9537
rect 46020 9571 46072 9580
rect 46020 9537 46029 9571
rect 46029 9537 46063 9571
rect 46063 9537 46072 9571
rect 46020 9528 46072 9537
rect 45560 9460 45612 9512
rect 46204 9460 46256 9512
rect 46848 9528 46900 9580
rect 48872 9571 48924 9580
rect 49240 9596 49292 9648
rect 50252 9639 50304 9648
rect 50252 9605 50261 9639
rect 50261 9605 50295 9639
rect 50295 9605 50304 9639
rect 50252 9596 50304 9605
rect 50896 9596 50948 9648
rect 51908 9639 51960 9648
rect 51908 9605 51917 9639
rect 51917 9605 51951 9639
rect 51951 9605 51960 9639
rect 51908 9596 51960 9605
rect 48872 9537 48911 9571
rect 48911 9537 48924 9571
rect 48872 9528 48924 9537
rect 48320 9460 48372 9512
rect 49792 9528 49844 9580
rect 50068 9528 50120 9580
rect 34612 9324 34664 9376
rect 35348 9324 35400 9376
rect 36176 9367 36228 9376
rect 36176 9333 36185 9367
rect 36185 9333 36219 9367
rect 36219 9333 36228 9367
rect 36176 9324 36228 9333
rect 36912 9324 36964 9376
rect 37648 9367 37700 9376
rect 37648 9333 37657 9367
rect 37657 9333 37691 9367
rect 37691 9333 37700 9367
rect 37648 9324 37700 9333
rect 38568 9324 38620 9376
rect 42432 9324 42484 9376
rect 42616 9367 42668 9376
rect 42616 9333 42625 9367
rect 42625 9333 42659 9367
rect 42659 9333 42668 9367
rect 42616 9324 42668 9333
rect 43720 9324 43772 9376
rect 46480 9392 46532 9444
rect 46940 9324 46992 9376
rect 48136 9392 48188 9444
rect 48964 9392 49016 9444
rect 52736 9596 52788 9648
rect 52920 9596 52972 9648
rect 52460 9528 52512 9580
rect 53288 9528 53340 9580
rect 52552 9460 52604 9512
rect 53472 9571 53524 9580
rect 53472 9537 53481 9571
rect 53481 9537 53515 9571
rect 53515 9537 53524 9571
rect 53472 9528 53524 9537
rect 53656 9528 53708 9580
rect 56048 9596 56100 9648
rect 56876 9596 56928 9648
rect 58072 9639 58124 9648
rect 58072 9605 58081 9639
rect 58081 9605 58115 9639
rect 58115 9605 58124 9639
rect 58072 9596 58124 9605
rect 56416 9571 56468 9580
rect 56416 9537 56425 9571
rect 56425 9537 56459 9571
rect 56459 9537 56468 9571
rect 56416 9528 56468 9537
rect 53748 9460 53800 9512
rect 54576 9460 54628 9512
rect 53012 9392 53064 9444
rect 55496 9435 55548 9444
rect 55496 9401 55505 9435
rect 55505 9401 55539 9435
rect 55539 9401 55548 9435
rect 55496 9392 55548 9401
rect 56876 9435 56928 9444
rect 56876 9401 56885 9435
rect 56885 9401 56919 9435
rect 56919 9401 56928 9435
rect 56876 9392 56928 9401
rect 49976 9324 50028 9376
rect 51080 9324 51132 9376
rect 54024 9324 54076 9376
rect 54852 9324 54904 9376
rect 56784 9324 56836 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 25964 9052 26016 9104
rect 27804 9052 27856 9104
rect 25688 8984 25740 9036
rect 28264 9052 28316 9104
rect 28908 9052 28960 9104
rect 29368 9052 29420 9104
rect 30288 9052 30340 9104
rect 30840 9120 30892 9172
rect 31576 9120 31628 9172
rect 32864 9120 32916 9172
rect 33048 9120 33100 9172
rect 33600 9120 33652 9172
rect 33876 9120 33928 9172
rect 34796 9120 34848 9172
rect 35072 9120 35124 9172
rect 35716 9120 35768 9172
rect 36452 9120 36504 9172
rect 31760 9052 31812 9104
rect 36728 9052 36780 9104
rect 37464 9120 37516 9172
rect 38384 9120 38436 9172
rect 38844 9163 38896 9172
rect 38844 9129 38853 9163
rect 38853 9129 38887 9163
rect 38887 9129 38896 9163
rect 38844 9120 38896 9129
rect 40684 9120 40736 9172
rect 46388 9120 46440 9172
rect 26056 8916 26108 8968
rect 26976 8916 27028 8968
rect 27620 8916 27672 8968
rect 27896 8959 27948 8968
rect 27896 8925 27905 8959
rect 27905 8925 27939 8959
rect 27939 8925 27948 8959
rect 27896 8916 27948 8925
rect 29828 8984 29880 9036
rect 30012 8984 30064 9036
rect 31576 8984 31628 9036
rect 35256 8984 35308 9036
rect 29000 8916 29052 8968
rect 29092 8916 29144 8968
rect 29644 8916 29696 8968
rect 30380 8959 30432 8968
rect 24032 8823 24084 8832
rect 24032 8789 24041 8823
rect 24041 8789 24075 8823
rect 24075 8789 24084 8823
rect 24032 8780 24084 8789
rect 25596 8780 25648 8832
rect 26516 8848 26568 8900
rect 26332 8780 26384 8832
rect 26792 8780 26844 8832
rect 27252 8848 27304 8900
rect 28448 8848 28500 8900
rect 29552 8848 29604 8900
rect 30380 8925 30389 8959
rect 30389 8925 30423 8959
rect 30423 8925 30432 8959
rect 30380 8916 30432 8925
rect 31392 8916 31444 8968
rect 32036 8848 32088 8900
rect 32312 8891 32364 8900
rect 30840 8780 30892 8832
rect 31392 8780 31444 8832
rect 31668 8780 31720 8832
rect 31852 8780 31904 8832
rect 32312 8857 32321 8891
rect 32321 8857 32355 8891
rect 32355 8857 32364 8891
rect 32312 8848 32364 8857
rect 32220 8780 32272 8832
rect 32956 8916 33008 8968
rect 33600 8959 33652 8968
rect 33600 8925 33609 8959
rect 33609 8925 33643 8959
rect 33643 8925 33652 8959
rect 33600 8916 33652 8925
rect 34152 8916 34204 8968
rect 34612 8916 34664 8968
rect 34796 8916 34848 8968
rect 35072 8959 35124 8968
rect 35072 8925 35081 8959
rect 35081 8925 35115 8959
rect 35115 8925 35124 8959
rect 35072 8916 35124 8925
rect 35348 8916 35400 8968
rect 36636 8984 36688 9036
rect 36912 8959 36964 8968
rect 36912 8925 36921 8959
rect 36921 8925 36955 8959
rect 36955 8925 36964 8959
rect 36912 8916 36964 8925
rect 35808 8848 35860 8900
rect 39580 8984 39632 9036
rect 37096 8959 37148 8968
rect 37096 8925 37105 8959
rect 37105 8925 37139 8959
rect 37139 8925 37148 8959
rect 37096 8916 37148 8925
rect 38936 8916 38988 8968
rect 40592 9052 40644 9104
rect 42524 9052 42576 9104
rect 42800 9052 42852 9104
rect 43536 9052 43588 9104
rect 45100 9052 45152 9104
rect 47032 9095 47084 9104
rect 47032 9061 47041 9095
rect 47041 9061 47075 9095
rect 47075 9061 47084 9095
rect 50252 9120 50304 9172
rect 50804 9163 50856 9172
rect 50804 9129 50813 9163
rect 50813 9129 50847 9163
rect 50847 9129 50856 9163
rect 50804 9120 50856 9129
rect 54208 9120 54260 9172
rect 55680 9120 55732 9172
rect 56600 9120 56652 9172
rect 47032 9052 47084 9061
rect 49608 9052 49660 9104
rect 49792 9052 49844 9104
rect 51356 9052 51408 9104
rect 51540 9052 51592 9104
rect 40408 8984 40460 9036
rect 41328 9027 41380 9036
rect 41328 8993 41337 9027
rect 41337 8993 41371 9027
rect 41371 8993 41380 9027
rect 41328 8984 41380 8993
rect 41052 8959 41104 8968
rect 41052 8925 41061 8959
rect 41061 8925 41095 8959
rect 41095 8925 41104 8959
rect 41052 8916 41104 8925
rect 41144 8959 41196 8968
rect 41144 8925 41153 8959
rect 41153 8925 41187 8959
rect 41187 8925 41196 8959
rect 41144 8916 41196 8925
rect 41788 8916 41840 8968
rect 43628 8984 43680 9036
rect 44916 8984 44968 9036
rect 45928 8984 45980 9036
rect 46020 8984 46072 9036
rect 42156 8959 42208 8968
rect 42156 8925 42166 8959
rect 42166 8925 42200 8959
rect 42200 8925 42208 8959
rect 42156 8916 42208 8925
rect 38384 8891 38436 8900
rect 38384 8857 38393 8891
rect 38393 8857 38427 8891
rect 38427 8857 38436 8891
rect 38384 8848 38436 8857
rect 39764 8848 39816 8900
rect 40408 8891 40460 8900
rect 40408 8857 40417 8891
rect 40417 8857 40451 8891
rect 40451 8857 40460 8891
rect 40408 8848 40460 8857
rect 43444 8848 43496 8900
rect 43628 8848 43680 8900
rect 44824 8916 44876 8968
rect 45284 8916 45336 8968
rect 45560 8848 45612 8900
rect 46112 8959 46164 8968
rect 46112 8925 46121 8959
rect 46121 8925 46155 8959
rect 46155 8925 46164 8959
rect 46112 8916 46164 8925
rect 46296 8959 46348 8968
rect 46296 8925 46305 8959
rect 46305 8925 46339 8959
rect 46339 8925 46348 8959
rect 46296 8916 46348 8925
rect 34336 8823 34388 8832
rect 34336 8789 34345 8823
rect 34345 8789 34379 8823
rect 34379 8789 34388 8823
rect 34336 8780 34388 8789
rect 34980 8823 35032 8832
rect 34980 8789 34989 8823
rect 34989 8789 35023 8823
rect 35023 8789 35032 8823
rect 34980 8780 35032 8789
rect 35992 8780 36044 8832
rect 37464 8780 37516 8832
rect 40132 8780 40184 8832
rect 43168 8780 43220 8832
rect 44088 8780 44140 8832
rect 44640 8780 44692 8832
rect 46204 8848 46256 8900
rect 46572 8780 46624 8832
rect 47216 8916 47268 8968
rect 48504 8916 48556 8968
rect 50068 8984 50120 9036
rect 49240 8916 49292 8968
rect 49976 8916 50028 8968
rect 52552 8984 52604 9036
rect 53932 9027 53984 9036
rect 53932 8993 53941 9027
rect 53941 8993 53975 9027
rect 53975 8993 53984 9027
rect 53932 8984 53984 8993
rect 54024 9027 54076 9036
rect 54024 8993 54033 9027
rect 54033 8993 54067 9027
rect 54067 8993 54076 9027
rect 54484 9052 54536 9104
rect 56324 9052 56376 9104
rect 54024 8984 54076 8993
rect 47584 8823 47636 8832
rect 47584 8789 47593 8823
rect 47593 8789 47627 8823
rect 47627 8789 47636 8823
rect 47584 8780 47636 8789
rect 47768 8780 47820 8832
rect 48136 8780 48188 8832
rect 49608 8848 49660 8900
rect 51724 8848 51776 8900
rect 52644 8916 52696 8968
rect 55404 8984 55456 9036
rect 48320 8780 48372 8832
rect 49148 8780 49200 8832
rect 50896 8780 50948 8832
rect 51172 8780 51224 8832
rect 52736 8848 52788 8900
rect 54392 8916 54444 8968
rect 56508 8916 56560 8968
rect 57336 8848 57388 8900
rect 53012 8780 53064 8832
rect 54576 8780 54628 8832
rect 56692 8823 56744 8832
rect 56692 8789 56701 8823
rect 56701 8789 56735 8823
rect 56735 8789 56744 8823
rect 56692 8780 56744 8789
rect 56876 8780 56928 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 25320 8576 25372 8628
rect 26700 8576 26752 8628
rect 28632 8576 28684 8628
rect 25596 8551 25648 8560
rect 25596 8517 25605 8551
rect 25605 8517 25639 8551
rect 25639 8517 25648 8551
rect 25596 8508 25648 8517
rect 25872 8508 25924 8560
rect 26608 8551 26660 8560
rect 26608 8517 26617 8551
rect 26617 8517 26651 8551
rect 26651 8517 26660 8551
rect 26608 8508 26660 8517
rect 25320 8483 25372 8492
rect 25320 8449 25329 8483
rect 25329 8449 25363 8483
rect 25363 8449 25372 8483
rect 25320 8440 25372 8449
rect 27160 8483 27212 8492
rect 27160 8449 27169 8483
rect 27169 8449 27203 8483
rect 27203 8449 27212 8483
rect 27160 8440 27212 8449
rect 28264 8508 28316 8560
rect 30196 8508 30248 8560
rect 28448 8440 28500 8492
rect 28632 8440 28684 8492
rect 29276 8440 29328 8492
rect 29552 8440 29604 8492
rect 30012 8440 30064 8492
rect 31300 8576 31352 8628
rect 37096 8576 37148 8628
rect 37556 8619 37608 8628
rect 37556 8585 37565 8619
rect 37565 8585 37599 8619
rect 37599 8585 37608 8619
rect 37556 8576 37608 8585
rect 38936 8619 38988 8628
rect 38936 8585 38945 8619
rect 38945 8585 38979 8619
rect 38979 8585 38988 8619
rect 38936 8576 38988 8585
rect 43996 8619 44048 8628
rect 43996 8585 44005 8619
rect 44005 8585 44039 8619
rect 44039 8585 44048 8619
rect 43996 8576 44048 8585
rect 46112 8576 46164 8628
rect 48320 8576 48372 8628
rect 49792 8576 49844 8628
rect 50712 8619 50764 8628
rect 50712 8585 50721 8619
rect 50721 8585 50755 8619
rect 50755 8585 50764 8619
rect 50712 8576 50764 8585
rect 51356 8576 51408 8628
rect 53012 8576 53064 8628
rect 53196 8576 53248 8628
rect 54024 8576 54076 8628
rect 54668 8619 54720 8628
rect 54668 8585 54677 8619
rect 54677 8585 54711 8619
rect 54711 8585 54720 8619
rect 54668 8576 54720 8585
rect 54852 8576 54904 8628
rect 55312 8576 55364 8628
rect 56692 8576 56744 8628
rect 30472 8508 30524 8560
rect 32496 8508 32548 8560
rect 32864 8508 32916 8560
rect 31392 8440 31444 8492
rect 31852 8440 31904 8492
rect 33232 8440 33284 8492
rect 33600 8440 33652 8492
rect 34980 8508 35032 8560
rect 35716 8508 35768 8560
rect 24032 8372 24084 8424
rect 26332 8372 26384 8424
rect 27436 8415 27488 8424
rect 27436 8381 27445 8415
rect 27445 8381 27479 8415
rect 27479 8381 27488 8415
rect 27436 8372 27488 8381
rect 30288 8372 30340 8424
rect 30472 8372 30524 8424
rect 30840 8372 30892 8424
rect 32772 8372 32824 8424
rect 32864 8415 32916 8424
rect 32864 8381 32873 8415
rect 32873 8381 32907 8415
rect 32907 8381 32916 8415
rect 32864 8372 32916 8381
rect 33692 8372 33744 8424
rect 34520 8440 34572 8492
rect 35256 8483 35308 8492
rect 35256 8449 35265 8483
rect 35265 8449 35299 8483
rect 35299 8449 35308 8483
rect 35440 8483 35492 8492
rect 35256 8440 35308 8449
rect 35440 8449 35449 8483
rect 35449 8449 35483 8483
rect 35483 8449 35492 8483
rect 35440 8440 35492 8449
rect 35624 8483 35676 8492
rect 35624 8449 35633 8483
rect 35633 8449 35667 8483
rect 35667 8449 35676 8483
rect 35624 8440 35676 8449
rect 35900 8440 35952 8492
rect 42984 8508 43036 8560
rect 46204 8551 46256 8560
rect 46204 8517 46213 8551
rect 46213 8517 46247 8551
rect 46247 8517 46256 8551
rect 46204 8508 46256 8517
rect 46572 8508 46624 8560
rect 36728 8483 36780 8492
rect 36728 8449 36737 8483
rect 36737 8449 36771 8483
rect 36771 8449 36780 8483
rect 36728 8440 36780 8449
rect 37740 8483 37792 8492
rect 37740 8449 37749 8483
rect 37749 8449 37783 8483
rect 37783 8449 37792 8483
rect 37740 8440 37792 8449
rect 38200 8440 38252 8492
rect 38568 8440 38620 8492
rect 39396 8483 39448 8492
rect 26424 8304 26476 8356
rect 28356 8304 28408 8356
rect 29184 8304 29236 8356
rect 30012 8304 30064 8356
rect 34152 8372 34204 8424
rect 34704 8372 34756 8424
rect 37280 8372 37332 8424
rect 38660 8372 38712 8424
rect 39396 8449 39405 8483
rect 39405 8449 39439 8483
rect 39439 8449 39448 8483
rect 39396 8440 39448 8449
rect 39580 8483 39632 8492
rect 39580 8449 39589 8483
rect 39589 8449 39623 8483
rect 39623 8449 39632 8483
rect 39580 8440 39632 8449
rect 40592 8483 40644 8492
rect 40592 8449 40601 8483
rect 40601 8449 40635 8483
rect 40635 8449 40644 8483
rect 40592 8440 40644 8449
rect 41788 8483 41840 8492
rect 41788 8449 41797 8483
rect 41797 8449 41831 8483
rect 41831 8449 41840 8483
rect 41788 8440 41840 8449
rect 42156 8440 42208 8492
rect 42984 8372 43036 8424
rect 43168 8415 43220 8424
rect 43168 8381 43177 8415
rect 43177 8381 43211 8415
rect 43211 8381 43220 8415
rect 43168 8372 43220 8381
rect 43536 8483 43588 8492
rect 43536 8449 43545 8483
rect 43545 8449 43579 8483
rect 43579 8449 43588 8483
rect 43536 8440 43588 8449
rect 44088 8440 44140 8492
rect 44916 8440 44968 8492
rect 45376 8440 45428 8492
rect 44456 8415 44508 8424
rect 34612 8304 34664 8356
rect 35532 8304 35584 8356
rect 40776 8347 40828 8356
rect 40776 8313 40785 8347
rect 40785 8313 40819 8347
rect 40819 8313 40828 8347
rect 40776 8304 40828 8313
rect 41604 8304 41656 8356
rect 44456 8381 44465 8415
rect 44465 8381 44499 8415
rect 44499 8381 44508 8415
rect 44456 8372 44508 8381
rect 44548 8415 44600 8424
rect 44548 8381 44557 8415
rect 44557 8381 44591 8415
rect 44591 8381 44600 8415
rect 44548 8372 44600 8381
rect 46020 8440 46072 8492
rect 46664 8440 46716 8492
rect 46848 8440 46900 8492
rect 45560 8372 45612 8424
rect 47584 8440 47636 8492
rect 48136 8440 48188 8492
rect 49608 8483 49660 8492
rect 49608 8449 49617 8483
rect 49617 8449 49651 8483
rect 49651 8449 49660 8483
rect 49608 8440 49660 8449
rect 50252 8508 50304 8560
rect 51448 8508 51500 8560
rect 54576 8508 54628 8560
rect 50068 8483 50120 8492
rect 50068 8449 50077 8483
rect 50077 8449 50111 8483
rect 50111 8449 50120 8483
rect 50068 8440 50120 8449
rect 48320 8415 48372 8424
rect 48320 8381 48329 8415
rect 48329 8381 48363 8415
rect 48363 8381 48372 8415
rect 48320 8372 48372 8381
rect 49792 8415 49844 8424
rect 49792 8381 49801 8415
rect 49801 8381 49835 8415
rect 49835 8381 49844 8415
rect 49792 8372 49844 8381
rect 46572 8304 46624 8356
rect 47124 8347 47176 8356
rect 47124 8313 47133 8347
rect 47133 8313 47167 8347
rect 47167 8313 47176 8347
rect 47124 8304 47176 8313
rect 2320 8236 2372 8288
rect 26884 8236 26936 8288
rect 29276 8236 29328 8288
rect 29920 8236 29972 8288
rect 33600 8279 33652 8288
rect 33600 8245 33609 8279
rect 33609 8245 33643 8279
rect 33643 8245 33652 8279
rect 33600 8236 33652 8245
rect 36176 8236 36228 8288
rect 37372 8236 37424 8288
rect 38844 8236 38896 8288
rect 40408 8279 40460 8288
rect 40408 8245 40417 8279
rect 40417 8245 40451 8279
rect 40451 8245 40460 8279
rect 40408 8236 40460 8245
rect 45284 8279 45336 8288
rect 45284 8245 45293 8279
rect 45293 8245 45327 8279
rect 45327 8245 45336 8279
rect 45284 8236 45336 8245
rect 46940 8236 46992 8288
rect 48136 8236 48188 8288
rect 49700 8236 49752 8288
rect 50160 8372 50212 8424
rect 50804 8372 50856 8424
rect 51448 8372 51500 8424
rect 51540 8372 51592 8424
rect 51908 8372 51960 8424
rect 52184 8440 52236 8492
rect 52920 8483 52972 8492
rect 52920 8449 52929 8483
rect 52929 8449 52963 8483
rect 52963 8449 52972 8483
rect 52920 8440 52972 8449
rect 50620 8304 50672 8356
rect 54852 8440 54904 8492
rect 54024 8372 54076 8424
rect 55496 8440 55548 8492
rect 56048 8440 56100 8492
rect 56416 8483 56468 8492
rect 56416 8449 56425 8483
rect 56425 8449 56459 8483
rect 56459 8449 56468 8483
rect 56416 8440 56468 8449
rect 57152 8440 57204 8492
rect 54300 8304 54352 8356
rect 55404 8347 55456 8356
rect 55404 8313 55413 8347
rect 55413 8313 55447 8347
rect 55447 8313 55456 8347
rect 55404 8304 55456 8313
rect 50896 8279 50948 8288
rect 50896 8245 50905 8279
rect 50905 8245 50939 8279
rect 50939 8245 50948 8279
rect 50896 8236 50948 8245
rect 50988 8236 51040 8288
rect 54392 8236 54444 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 25320 8032 25372 8084
rect 27436 8075 27488 8084
rect 27436 8041 27445 8075
rect 27445 8041 27479 8075
rect 27479 8041 27488 8075
rect 27436 8032 27488 8041
rect 27804 8032 27856 8084
rect 32956 8032 33008 8084
rect 33692 8032 33744 8084
rect 34612 8032 34664 8084
rect 35440 8032 35492 8084
rect 35624 8032 35676 8084
rect 35992 8075 36044 8084
rect 35992 8041 36001 8075
rect 36001 8041 36035 8075
rect 36035 8041 36044 8075
rect 35992 8032 36044 8041
rect 36268 8032 36320 8084
rect 37740 8032 37792 8084
rect 38660 8032 38712 8084
rect 39028 8032 39080 8084
rect 40500 8032 40552 8084
rect 40960 8075 41012 8084
rect 40960 8041 40969 8075
rect 40969 8041 41003 8075
rect 41003 8041 41012 8075
rect 40960 8032 41012 8041
rect 41328 8032 41380 8084
rect 42524 8032 42576 8084
rect 46480 8032 46532 8084
rect 46572 8032 46624 8084
rect 47860 8032 47912 8084
rect 48412 8032 48464 8084
rect 49884 8032 49936 8084
rect 50804 8032 50856 8084
rect 51816 8075 51868 8084
rect 25780 8007 25832 8016
rect 25780 7973 25789 8007
rect 25789 7973 25823 8007
rect 25823 7973 25832 8007
rect 25780 7964 25832 7973
rect 27252 7964 27304 8016
rect 28816 7964 28868 8016
rect 32772 7964 32824 8016
rect 33140 7964 33192 8016
rect 38936 8007 38988 8016
rect 25228 7871 25280 7880
rect 25228 7837 25237 7871
rect 25237 7837 25271 7871
rect 25271 7837 25280 7871
rect 25412 7871 25464 7880
rect 25228 7828 25280 7837
rect 25412 7837 25430 7871
rect 25430 7837 25464 7871
rect 25412 7828 25464 7837
rect 26516 7896 26568 7948
rect 26792 7896 26844 7948
rect 26884 7896 26936 7948
rect 35164 7939 35216 7948
rect 26976 7871 27028 7880
rect 26976 7837 26985 7871
rect 26985 7837 27019 7871
rect 27019 7837 27028 7871
rect 26976 7828 27028 7837
rect 28540 7871 28592 7880
rect 28540 7837 28549 7871
rect 28549 7837 28583 7871
rect 28583 7837 28592 7871
rect 28540 7828 28592 7837
rect 29092 7828 29144 7880
rect 29552 7828 29604 7880
rect 29828 7871 29880 7880
rect 29828 7837 29837 7871
rect 29837 7837 29871 7871
rect 29871 7837 29880 7871
rect 29828 7828 29880 7837
rect 31484 7828 31536 7880
rect 31760 7871 31812 7880
rect 31760 7837 31769 7871
rect 31769 7837 31803 7871
rect 31803 7837 31812 7871
rect 31760 7828 31812 7837
rect 32128 7871 32180 7880
rect 32128 7837 32137 7871
rect 32137 7837 32171 7871
rect 32171 7837 32180 7871
rect 32128 7828 32180 7837
rect 32496 7828 32548 7880
rect 33140 7871 33192 7880
rect 33140 7837 33149 7871
rect 33149 7837 33183 7871
rect 33183 7837 33192 7871
rect 33140 7828 33192 7837
rect 27528 7760 27580 7812
rect 28908 7760 28960 7812
rect 30288 7760 30340 7812
rect 28264 7692 28316 7744
rect 29000 7692 29052 7744
rect 29828 7692 29880 7744
rect 30472 7692 30524 7744
rect 30656 7735 30708 7744
rect 30656 7701 30665 7735
rect 30665 7701 30699 7735
rect 30699 7701 30708 7735
rect 30656 7692 30708 7701
rect 31116 7692 31168 7744
rect 32312 7760 32364 7812
rect 33600 7828 33652 7880
rect 34060 7871 34112 7880
rect 34060 7837 34069 7871
rect 34069 7837 34103 7871
rect 34103 7837 34112 7871
rect 34060 7828 34112 7837
rect 35164 7905 35173 7939
rect 35173 7905 35207 7939
rect 35207 7905 35216 7939
rect 35164 7896 35216 7905
rect 35900 7828 35952 7880
rect 36176 7871 36228 7880
rect 36176 7837 36185 7871
rect 36185 7837 36219 7871
rect 36219 7837 36228 7871
rect 36176 7828 36228 7837
rect 36728 7871 36780 7880
rect 36728 7837 36737 7871
rect 36737 7837 36771 7871
rect 36771 7837 36780 7871
rect 36728 7828 36780 7837
rect 37648 7828 37700 7880
rect 38016 7871 38068 7880
rect 38016 7837 38025 7871
rect 38025 7837 38059 7871
rect 38059 7837 38068 7871
rect 38016 7828 38068 7837
rect 38936 7973 38945 8007
rect 38945 7973 38979 8007
rect 38979 7973 38988 8007
rect 38936 7964 38988 7973
rect 39396 7964 39448 8016
rect 40224 7964 40276 8016
rect 42800 8007 42852 8016
rect 42800 7973 42809 8007
rect 42809 7973 42843 8007
rect 42843 7973 42852 8007
rect 42800 7964 42852 7973
rect 46388 7964 46440 8016
rect 51172 7964 51224 8016
rect 51356 7964 51408 8016
rect 51816 8041 51825 8075
rect 51825 8041 51859 8075
rect 51859 8041 51868 8075
rect 51816 8032 51868 8041
rect 52092 8032 52144 8084
rect 39580 7896 39632 7948
rect 42156 7896 42208 7948
rect 42708 7896 42760 7948
rect 41420 7828 41472 7880
rect 44088 7896 44140 7948
rect 46756 7896 46808 7948
rect 36544 7760 36596 7812
rect 41604 7760 41656 7812
rect 38200 7735 38252 7744
rect 38200 7701 38209 7735
rect 38209 7701 38243 7735
rect 38243 7701 38252 7735
rect 38200 7692 38252 7701
rect 41512 7735 41564 7744
rect 41512 7701 41521 7735
rect 41521 7701 41555 7735
rect 41555 7701 41564 7735
rect 41512 7692 41564 7701
rect 43260 7692 43312 7744
rect 44272 7828 44324 7880
rect 44456 7828 44508 7880
rect 46572 7871 46624 7880
rect 46572 7837 46581 7871
rect 46581 7837 46615 7871
rect 46615 7837 46624 7871
rect 46572 7828 46624 7837
rect 47584 7896 47636 7948
rect 44548 7760 44600 7812
rect 44088 7692 44140 7744
rect 45836 7692 45888 7744
rect 46296 7692 46348 7744
rect 46480 7692 46532 7744
rect 47676 7871 47728 7880
rect 47676 7837 47685 7871
rect 47685 7837 47719 7871
rect 47719 7837 47728 7871
rect 47676 7828 47728 7837
rect 47860 7871 47912 7880
rect 47860 7837 47869 7871
rect 47869 7837 47903 7871
rect 47903 7837 47912 7871
rect 47860 7828 47912 7837
rect 48136 7828 48188 7880
rect 49792 7896 49844 7948
rect 50068 7896 50120 7948
rect 50988 7896 51040 7948
rect 49332 7871 49384 7880
rect 49332 7837 49341 7871
rect 49341 7837 49375 7871
rect 49375 7837 49384 7871
rect 49332 7828 49384 7837
rect 49516 7871 49568 7880
rect 49516 7837 49525 7871
rect 49525 7837 49559 7871
rect 49559 7837 49568 7871
rect 49516 7828 49568 7837
rect 51908 7896 51960 7948
rect 48228 7760 48280 7812
rect 51540 7871 51592 7880
rect 49884 7760 49936 7812
rect 51540 7837 51549 7871
rect 51549 7837 51583 7871
rect 51583 7837 51592 7871
rect 51540 7828 51592 7837
rect 52000 7828 52052 7880
rect 51448 7760 51500 7812
rect 52276 7964 52328 8016
rect 53472 7896 53524 7948
rect 53012 7871 53064 7880
rect 53012 7837 53021 7871
rect 53021 7837 53055 7871
rect 53055 7837 53064 7871
rect 53012 7828 53064 7837
rect 53288 7828 53340 7880
rect 53656 7760 53708 7812
rect 54116 7828 54168 7880
rect 54392 7871 54444 7880
rect 54392 7837 54401 7871
rect 54401 7837 54435 7871
rect 54435 7837 54444 7871
rect 54392 7828 54444 7837
rect 56048 8032 56100 8084
rect 57428 8075 57480 8084
rect 57428 8041 57437 8075
rect 57437 8041 57471 8075
rect 57471 8041 57480 8075
rect 57428 8032 57480 8041
rect 54760 7964 54812 8016
rect 55128 7964 55180 8016
rect 55864 8007 55916 8016
rect 55864 7973 55873 8007
rect 55873 7973 55907 8007
rect 55907 7973 55916 8007
rect 55864 7964 55916 7973
rect 54852 7896 54904 7948
rect 56140 7896 56192 7948
rect 54760 7828 54812 7880
rect 55864 7828 55916 7880
rect 56784 7828 56836 7880
rect 49792 7692 49844 7744
rect 51080 7692 51132 7744
rect 51632 7692 51684 7744
rect 52644 7692 52696 7744
rect 55680 7692 55732 7744
rect 57980 7735 58032 7744
rect 57980 7701 57989 7735
rect 57989 7701 58023 7735
rect 58023 7701 58032 7735
rect 57980 7692 58032 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 23848 7420 23900 7472
rect 25412 7420 25464 7472
rect 25872 7488 25924 7540
rect 27068 7488 27120 7540
rect 26976 7420 27028 7472
rect 24952 7395 25004 7404
rect 24952 7361 24961 7395
rect 24961 7361 24995 7395
rect 24995 7361 25004 7395
rect 24952 7352 25004 7361
rect 25964 7395 26016 7404
rect 25964 7361 25973 7395
rect 25973 7361 26007 7395
rect 26007 7361 26016 7395
rect 25964 7352 26016 7361
rect 26240 7395 26292 7404
rect 26240 7361 26249 7395
rect 26249 7361 26283 7395
rect 26283 7361 26292 7395
rect 26240 7352 26292 7361
rect 26332 7395 26384 7404
rect 26332 7361 26341 7395
rect 26341 7361 26375 7395
rect 26375 7361 26384 7395
rect 26332 7352 26384 7361
rect 27620 7395 27672 7404
rect 27620 7361 27629 7395
rect 27629 7361 27663 7395
rect 27663 7361 27672 7395
rect 27620 7352 27672 7361
rect 28724 7420 28776 7472
rect 31576 7488 31628 7540
rect 32496 7488 32548 7540
rect 35348 7488 35400 7540
rect 35624 7531 35676 7540
rect 35624 7497 35633 7531
rect 35633 7497 35667 7531
rect 35667 7497 35676 7531
rect 35624 7488 35676 7497
rect 36636 7488 36688 7540
rect 29092 7352 29144 7404
rect 29460 7395 29512 7404
rect 29460 7361 29469 7395
rect 29469 7361 29503 7395
rect 29503 7361 29512 7395
rect 29460 7352 29512 7361
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 30472 7395 30524 7404
rect 30472 7361 30481 7395
rect 30481 7361 30515 7395
rect 30515 7361 30524 7395
rect 30472 7352 30524 7361
rect 31300 7352 31352 7404
rect 31484 7352 31536 7404
rect 32036 7352 32088 7404
rect 32864 7420 32916 7472
rect 35716 7420 35768 7472
rect 38936 7488 38988 7540
rect 40408 7488 40460 7540
rect 42800 7488 42852 7540
rect 43352 7488 43404 7540
rect 44456 7488 44508 7540
rect 45744 7488 45796 7540
rect 37464 7463 37516 7472
rect 37464 7429 37473 7463
rect 37473 7429 37507 7463
rect 37507 7429 37516 7463
rect 37464 7420 37516 7429
rect 38016 7420 38068 7472
rect 39580 7420 39632 7472
rect 33600 7352 33652 7404
rect 33784 7395 33836 7404
rect 33784 7361 33793 7395
rect 33793 7361 33827 7395
rect 33827 7361 33836 7395
rect 33784 7352 33836 7361
rect 33968 7395 34020 7404
rect 33968 7361 33977 7395
rect 33977 7361 34011 7395
rect 34011 7361 34020 7395
rect 33968 7352 34020 7361
rect 26700 7284 26752 7336
rect 26976 7284 27028 7336
rect 27896 7284 27948 7336
rect 27988 7284 28040 7336
rect 28448 7284 28500 7336
rect 28908 7284 28960 7336
rect 30288 7284 30340 7336
rect 32496 7327 32548 7336
rect 27436 7259 27488 7268
rect 27436 7225 27445 7259
rect 27445 7225 27479 7259
rect 27479 7225 27488 7259
rect 27436 7216 27488 7225
rect 25136 7148 25188 7200
rect 26240 7148 26292 7200
rect 30104 7216 30156 7268
rect 30196 7216 30248 7268
rect 32496 7293 32505 7327
rect 32505 7293 32539 7327
rect 32539 7293 32548 7327
rect 32496 7284 32548 7293
rect 32680 7327 32732 7336
rect 32680 7293 32689 7327
rect 32689 7293 32723 7327
rect 32723 7293 32732 7327
rect 32680 7284 32732 7293
rect 32772 7284 32824 7336
rect 30840 7216 30892 7268
rect 33692 7216 33744 7268
rect 27712 7148 27764 7200
rect 31668 7148 31720 7200
rect 33232 7148 33284 7200
rect 33508 7191 33560 7200
rect 33508 7157 33517 7191
rect 33517 7157 33551 7191
rect 33551 7157 33560 7191
rect 33508 7148 33560 7157
rect 35348 7284 35400 7336
rect 35900 7352 35952 7404
rect 36636 7395 36688 7404
rect 36636 7361 36645 7395
rect 36645 7361 36679 7395
rect 36679 7361 36688 7395
rect 36636 7352 36688 7361
rect 37004 7284 37056 7336
rect 38292 7395 38344 7404
rect 38292 7361 38301 7395
rect 38301 7361 38335 7395
rect 38335 7361 38344 7395
rect 38292 7352 38344 7361
rect 38660 7352 38712 7404
rect 40684 7420 40736 7472
rect 43996 7463 44048 7472
rect 43996 7429 44005 7463
rect 44005 7429 44039 7463
rect 44039 7429 44048 7463
rect 43996 7420 44048 7429
rect 46296 7463 46348 7472
rect 46296 7429 46305 7463
rect 46305 7429 46339 7463
rect 46339 7429 46348 7463
rect 46296 7420 46348 7429
rect 46388 7463 46440 7472
rect 46388 7429 46397 7463
rect 46397 7429 46431 7463
rect 46431 7429 46440 7463
rect 46388 7420 46440 7429
rect 46940 7420 46992 7472
rect 48136 7488 48188 7540
rect 40960 7395 41012 7404
rect 38016 7327 38068 7336
rect 38016 7293 38025 7327
rect 38025 7293 38059 7327
rect 38059 7293 38068 7327
rect 38016 7284 38068 7293
rect 39396 7284 39448 7336
rect 40960 7361 40969 7395
rect 40969 7361 41003 7395
rect 41003 7361 41012 7395
rect 40960 7352 41012 7361
rect 42892 7395 42944 7404
rect 42892 7361 42901 7395
rect 42901 7361 42935 7395
rect 42935 7361 42944 7395
rect 42892 7352 42944 7361
rect 42984 7395 43036 7404
rect 42984 7361 42993 7395
rect 42993 7361 43027 7395
rect 43027 7361 43036 7395
rect 42984 7352 43036 7361
rect 43168 7352 43220 7404
rect 44088 7352 44140 7404
rect 44180 7352 44232 7404
rect 44916 7352 44968 7404
rect 46204 7395 46256 7404
rect 46204 7361 46213 7395
rect 46213 7361 46247 7395
rect 46247 7361 46256 7395
rect 46204 7352 46256 7361
rect 47216 7352 47268 7404
rect 47584 7352 47636 7404
rect 34152 7216 34204 7268
rect 35532 7259 35584 7268
rect 35532 7225 35541 7259
rect 35541 7225 35575 7259
rect 35575 7225 35584 7259
rect 35532 7216 35584 7225
rect 37096 7216 37148 7268
rect 42524 7284 42576 7336
rect 43444 7284 43496 7336
rect 46388 7284 46440 7336
rect 48412 7420 48464 7472
rect 50068 7488 50120 7540
rect 51540 7488 51592 7540
rect 52552 7488 52604 7540
rect 52736 7488 52788 7540
rect 51264 7420 51316 7472
rect 53932 7488 53984 7540
rect 54208 7531 54260 7540
rect 54208 7497 54217 7531
rect 54217 7497 54251 7531
rect 54251 7497 54260 7531
rect 54208 7488 54260 7497
rect 56784 7488 56836 7540
rect 48596 7352 48648 7404
rect 48872 7352 48924 7404
rect 48964 7352 49016 7404
rect 49792 7395 49844 7404
rect 49792 7361 49801 7395
rect 49801 7361 49835 7395
rect 49835 7361 49844 7395
rect 49792 7352 49844 7361
rect 51356 7352 51408 7404
rect 52184 7352 52236 7404
rect 49608 7327 49660 7336
rect 37464 7148 37516 7200
rect 38568 7148 38620 7200
rect 40500 7216 40552 7268
rect 40684 7216 40736 7268
rect 41052 7148 41104 7200
rect 41972 7148 42024 7200
rect 44272 7216 44324 7268
rect 47860 7216 47912 7268
rect 49332 7216 49384 7268
rect 49608 7293 49617 7327
rect 49617 7293 49651 7327
rect 49651 7293 49660 7327
rect 49608 7284 49660 7293
rect 49884 7327 49936 7336
rect 49884 7293 49893 7327
rect 49893 7293 49927 7327
rect 49927 7293 49936 7327
rect 49884 7284 49936 7293
rect 51080 7327 51132 7336
rect 51080 7293 51089 7327
rect 51089 7293 51123 7327
rect 51123 7293 51132 7327
rect 52920 7395 52972 7404
rect 52920 7361 52929 7395
rect 52929 7361 52963 7395
rect 52963 7361 52972 7395
rect 52920 7352 52972 7361
rect 53472 7352 53524 7404
rect 54116 7420 54168 7472
rect 56140 7420 56192 7472
rect 53932 7352 53984 7404
rect 54484 7395 54536 7404
rect 54484 7361 54493 7395
rect 54493 7361 54527 7395
rect 54527 7361 54536 7395
rect 54484 7352 54536 7361
rect 54668 7395 54720 7404
rect 54668 7361 54677 7395
rect 54677 7361 54711 7395
rect 54711 7361 54720 7395
rect 54668 7352 54720 7361
rect 54852 7395 54904 7404
rect 54852 7361 54861 7395
rect 54861 7361 54895 7395
rect 54895 7361 54904 7395
rect 58072 7395 58124 7404
rect 54852 7352 54904 7361
rect 58072 7361 58081 7395
rect 58081 7361 58115 7395
rect 58115 7361 58124 7395
rect 58072 7352 58124 7361
rect 51080 7284 51132 7293
rect 44364 7191 44416 7200
rect 44364 7157 44373 7191
rect 44373 7157 44407 7191
rect 44407 7157 44416 7191
rect 44364 7148 44416 7157
rect 45284 7148 45336 7200
rect 47032 7148 47084 7200
rect 49424 7191 49476 7200
rect 49424 7157 49433 7191
rect 49433 7157 49467 7191
rect 49467 7157 49476 7191
rect 49424 7148 49476 7157
rect 49792 7148 49844 7200
rect 53288 7284 53340 7336
rect 54300 7284 54352 7336
rect 56968 7216 57020 7268
rect 51724 7148 51776 7200
rect 52736 7148 52788 7200
rect 53380 7191 53432 7200
rect 53380 7157 53389 7191
rect 53389 7157 53423 7191
rect 53423 7157 53432 7191
rect 53380 7148 53432 7157
rect 53656 7148 53708 7200
rect 54760 7191 54812 7200
rect 54760 7157 54769 7191
rect 54769 7157 54803 7191
rect 54803 7157 54812 7191
rect 54760 7148 54812 7157
rect 55496 7191 55548 7200
rect 55496 7157 55505 7191
rect 55505 7157 55539 7191
rect 55539 7157 55548 7191
rect 55496 7148 55548 7157
rect 55680 7148 55732 7200
rect 56324 7148 56376 7200
rect 57888 7148 57940 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 27436 6944 27488 6996
rect 27620 6944 27672 6996
rect 28356 6944 28408 6996
rect 30840 6944 30892 6996
rect 34060 6944 34112 6996
rect 34152 6944 34204 6996
rect 34796 6944 34848 6996
rect 35440 6944 35492 6996
rect 38660 6944 38712 6996
rect 41144 6944 41196 6996
rect 43720 6944 43772 6996
rect 45560 6944 45612 6996
rect 45744 6944 45796 6996
rect 46940 6944 46992 6996
rect 47216 6987 47268 6996
rect 47216 6953 47225 6987
rect 47225 6953 47259 6987
rect 47259 6953 47268 6987
rect 47216 6944 47268 6953
rect 48228 6944 48280 6996
rect 48596 6944 48648 6996
rect 49424 6944 49476 6996
rect 24308 6876 24360 6928
rect 27068 6876 27120 6928
rect 27252 6876 27304 6928
rect 28816 6876 28868 6928
rect 29644 6876 29696 6928
rect 31116 6876 31168 6928
rect 25044 6783 25096 6792
rect 25044 6749 25053 6783
rect 25053 6749 25087 6783
rect 25087 6749 25096 6783
rect 25044 6740 25096 6749
rect 25136 6783 25188 6792
rect 25136 6749 25146 6783
rect 25146 6749 25180 6783
rect 25180 6749 25188 6783
rect 25136 6740 25188 6749
rect 25872 6740 25924 6792
rect 24952 6672 25004 6724
rect 26332 6740 26384 6792
rect 26700 6740 26752 6792
rect 26148 6672 26200 6724
rect 26792 6715 26844 6724
rect 25504 6604 25556 6656
rect 26792 6681 26801 6715
rect 26801 6681 26835 6715
rect 26835 6681 26844 6715
rect 26792 6672 26844 6681
rect 27436 6740 27488 6792
rect 27528 6783 27580 6792
rect 27528 6749 27537 6783
rect 27537 6749 27571 6783
rect 27571 6749 27580 6783
rect 27528 6740 27580 6749
rect 27252 6715 27304 6724
rect 27252 6681 27261 6715
rect 27261 6681 27295 6715
rect 27295 6681 27304 6715
rect 27252 6672 27304 6681
rect 28080 6808 28132 6860
rect 28540 6808 28592 6860
rect 29828 6851 29880 6860
rect 29828 6817 29837 6851
rect 29837 6817 29871 6851
rect 29871 6817 29880 6851
rect 29828 6808 29880 6817
rect 30196 6808 30248 6860
rect 31392 6808 31444 6860
rect 33600 6876 33652 6928
rect 34704 6876 34756 6928
rect 35624 6876 35676 6928
rect 34060 6808 34112 6860
rect 28356 6783 28408 6792
rect 28356 6749 28365 6783
rect 28365 6749 28399 6783
rect 28399 6749 28408 6783
rect 28356 6740 28408 6749
rect 28448 6740 28500 6792
rect 27804 6672 27856 6724
rect 29644 6740 29696 6792
rect 30380 6672 30432 6724
rect 29920 6604 29972 6656
rect 30564 6740 30616 6792
rect 31024 6783 31076 6792
rect 31024 6749 31033 6783
rect 31033 6749 31067 6783
rect 31067 6749 31076 6783
rect 31024 6740 31076 6749
rect 31116 6740 31168 6792
rect 31852 6783 31904 6792
rect 31852 6749 31861 6783
rect 31861 6749 31895 6783
rect 31895 6749 31904 6783
rect 31852 6740 31904 6749
rect 32128 6740 32180 6792
rect 32680 6783 32732 6792
rect 32680 6749 32690 6783
rect 32690 6749 32724 6783
rect 32724 6749 32732 6783
rect 32680 6740 32732 6749
rect 33508 6740 33560 6792
rect 33600 6740 33652 6792
rect 33876 6740 33928 6792
rect 31668 6604 31720 6656
rect 32496 6647 32548 6656
rect 32496 6613 32505 6647
rect 32505 6613 32539 6647
rect 32539 6613 32548 6647
rect 32496 6604 32548 6613
rect 33140 6672 33192 6724
rect 34244 6808 34296 6860
rect 35716 6808 35768 6860
rect 35900 6740 35952 6792
rect 36084 6783 36136 6792
rect 36084 6749 36093 6783
rect 36093 6749 36127 6783
rect 36127 6749 36136 6783
rect 36084 6740 36136 6749
rect 36176 6740 36228 6792
rect 38292 6876 38344 6928
rect 41604 6876 41656 6928
rect 43628 6876 43680 6928
rect 46572 6876 46624 6928
rect 46664 6876 46716 6928
rect 50804 6944 50856 6996
rect 37188 6808 37240 6860
rect 37648 6740 37700 6792
rect 38016 6783 38068 6792
rect 38016 6749 38025 6783
rect 38025 6749 38059 6783
rect 38059 6749 38068 6783
rect 38016 6740 38068 6749
rect 39488 6783 39540 6792
rect 39488 6749 39497 6783
rect 39497 6749 39531 6783
rect 39531 6749 39540 6783
rect 39488 6740 39540 6749
rect 40224 6783 40276 6792
rect 40224 6749 40233 6783
rect 40233 6749 40267 6783
rect 40267 6749 40276 6783
rect 40224 6740 40276 6749
rect 40500 6740 40552 6792
rect 41972 6808 42024 6860
rect 42524 6851 42576 6860
rect 42524 6817 42533 6851
rect 42533 6817 42567 6851
rect 42567 6817 42576 6851
rect 42524 6808 42576 6817
rect 36728 6672 36780 6724
rect 37740 6672 37792 6724
rect 41420 6783 41472 6792
rect 41420 6749 41429 6783
rect 41429 6749 41463 6783
rect 41463 6749 41472 6783
rect 41420 6740 41472 6749
rect 42892 6808 42944 6860
rect 45376 6808 45428 6860
rect 46756 6808 46808 6860
rect 47400 6851 47452 6860
rect 47400 6817 47409 6851
rect 47409 6817 47443 6851
rect 47443 6817 47452 6851
rect 47400 6808 47452 6817
rect 42984 6672 43036 6724
rect 43904 6715 43956 6724
rect 39120 6604 39172 6656
rect 39304 6647 39356 6656
rect 39304 6613 39313 6647
rect 39313 6613 39347 6647
rect 39347 6613 39356 6647
rect 39304 6604 39356 6613
rect 40408 6647 40460 6656
rect 40408 6613 40417 6647
rect 40417 6613 40451 6647
rect 40451 6613 40460 6647
rect 40408 6604 40460 6613
rect 41420 6604 41472 6656
rect 43904 6681 43913 6715
rect 43913 6681 43947 6715
rect 43947 6681 43956 6715
rect 43904 6672 43956 6681
rect 44364 6672 44416 6724
rect 45284 6672 45336 6724
rect 45744 6715 45796 6724
rect 45744 6681 45753 6715
rect 45753 6681 45787 6715
rect 45787 6681 45796 6715
rect 47308 6783 47360 6792
rect 47308 6749 47317 6783
rect 47317 6749 47351 6783
rect 47351 6749 47360 6783
rect 47584 6783 47636 6792
rect 47308 6740 47360 6749
rect 47584 6749 47593 6783
rect 47593 6749 47627 6783
rect 47627 6749 47636 6783
rect 47584 6740 47636 6749
rect 47676 6783 47728 6792
rect 47676 6749 47685 6783
rect 47685 6749 47719 6783
rect 47719 6749 47728 6783
rect 47676 6740 47728 6749
rect 48044 6740 48096 6792
rect 50160 6876 50212 6928
rect 51264 6876 51316 6928
rect 49056 6851 49108 6860
rect 49056 6817 49065 6851
rect 49065 6817 49099 6851
rect 49099 6817 49108 6851
rect 49056 6808 49108 6817
rect 49792 6808 49844 6860
rect 52920 6944 52972 6996
rect 56324 6987 56376 6996
rect 52828 6876 52880 6928
rect 56324 6953 56333 6987
rect 56333 6953 56367 6987
rect 56367 6953 56376 6987
rect 56324 6944 56376 6953
rect 58072 6987 58124 6996
rect 58072 6953 58081 6987
rect 58081 6953 58115 6987
rect 58115 6953 58124 6987
rect 58072 6944 58124 6953
rect 54668 6919 54720 6928
rect 54668 6885 54677 6919
rect 54677 6885 54711 6919
rect 54711 6885 54720 6919
rect 54668 6876 54720 6885
rect 49332 6783 49384 6792
rect 49332 6749 49341 6783
rect 49341 6749 49375 6783
rect 49375 6749 49384 6783
rect 49332 6740 49384 6749
rect 49884 6740 49936 6792
rect 50344 6783 50396 6792
rect 50344 6749 50353 6783
rect 50353 6749 50387 6783
rect 50387 6749 50396 6783
rect 50344 6740 50396 6749
rect 50804 6740 50856 6792
rect 51724 6783 51776 6792
rect 51724 6749 51733 6783
rect 51733 6749 51767 6783
rect 51767 6749 51776 6783
rect 51724 6740 51776 6749
rect 51908 6783 51960 6792
rect 51908 6749 51917 6783
rect 51917 6749 51951 6783
rect 51951 6749 51960 6783
rect 51908 6740 51960 6749
rect 45744 6672 45796 6681
rect 48688 6672 48740 6724
rect 52460 6808 52512 6860
rect 55220 6808 55272 6860
rect 56232 6808 56284 6860
rect 57336 6808 57388 6860
rect 52276 6740 52328 6792
rect 54760 6740 54812 6792
rect 45928 6604 45980 6656
rect 46296 6604 46348 6656
rect 47400 6604 47452 6656
rect 52460 6672 52512 6724
rect 53288 6715 53340 6724
rect 52552 6604 52604 6656
rect 52736 6647 52788 6656
rect 52736 6613 52745 6647
rect 52745 6613 52779 6647
rect 52779 6613 52788 6647
rect 52736 6604 52788 6613
rect 53288 6681 53297 6715
rect 53297 6681 53331 6715
rect 53331 6681 53340 6715
rect 53288 6672 53340 6681
rect 54852 6715 54904 6724
rect 54852 6681 54861 6715
rect 54861 6681 54895 6715
rect 54895 6681 54904 6715
rect 54852 6672 54904 6681
rect 55036 6672 55088 6724
rect 58532 6740 58584 6792
rect 54116 6604 54168 6656
rect 54208 6604 54260 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 24124 6443 24176 6452
rect 24124 6409 24133 6443
rect 24133 6409 24167 6443
rect 24167 6409 24176 6443
rect 24124 6400 24176 6409
rect 25228 6400 25280 6452
rect 29000 6443 29052 6452
rect 29000 6409 29009 6443
rect 29009 6409 29043 6443
rect 29043 6409 29052 6443
rect 29000 6400 29052 6409
rect 29644 6443 29696 6452
rect 29644 6409 29653 6443
rect 29653 6409 29687 6443
rect 29687 6409 29696 6443
rect 29644 6400 29696 6409
rect 25412 6332 25464 6384
rect 28080 6332 28132 6384
rect 28356 6332 28408 6384
rect 25320 6307 25372 6316
rect 25320 6273 25329 6307
rect 25329 6273 25363 6307
rect 25363 6273 25372 6307
rect 25320 6264 25372 6273
rect 26056 6307 26108 6316
rect 25780 6196 25832 6248
rect 26056 6273 26065 6307
rect 26065 6273 26099 6307
rect 26099 6273 26108 6307
rect 26056 6264 26108 6273
rect 29828 6332 29880 6384
rect 26332 6196 26384 6248
rect 26700 6196 26752 6248
rect 27436 6196 27488 6248
rect 28356 6196 28408 6248
rect 30748 6332 30800 6384
rect 30932 6400 30984 6452
rect 32128 6400 32180 6452
rect 30564 6264 30616 6316
rect 31484 6332 31536 6384
rect 32588 6400 32640 6452
rect 34060 6400 34112 6452
rect 39856 6400 39908 6452
rect 32680 6332 32732 6384
rect 33140 6332 33192 6384
rect 33508 6332 33560 6384
rect 31300 6264 31352 6316
rect 31392 6264 31444 6316
rect 33692 6307 33744 6316
rect 33692 6273 33701 6307
rect 33701 6273 33735 6307
rect 33735 6273 33744 6307
rect 33692 6264 33744 6273
rect 34244 6264 34296 6316
rect 34612 6332 34664 6384
rect 36452 6375 36504 6384
rect 35716 6264 35768 6316
rect 36452 6341 36461 6375
rect 36461 6341 36495 6375
rect 36495 6341 36504 6375
rect 36452 6332 36504 6341
rect 38016 6332 38068 6384
rect 38200 6332 38252 6384
rect 38660 6332 38712 6384
rect 36360 6264 36412 6316
rect 36912 6307 36964 6316
rect 36912 6273 36921 6307
rect 36921 6273 36955 6307
rect 36955 6273 36964 6307
rect 36912 6264 36964 6273
rect 37096 6264 37148 6316
rect 38108 6264 38160 6316
rect 38844 6375 38896 6384
rect 38844 6341 38857 6375
rect 38857 6341 38891 6375
rect 38891 6341 38896 6375
rect 38844 6332 38896 6341
rect 38936 6307 38988 6316
rect 38936 6273 38945 6307
rect 38945 6273 38979 6307
rect 38979 6273 38988 6307
rect 38936 6264 38988 6273
rect 39120 6307 39172 6316
rect 39120 6273 39129 6307
rect 39129 6273 39163 6307
rect 39163 6273 39172 6307
rect 39856 6307 39908 6316
rect 39120 6264 39172 6273
rect 30380 6196 30432 6248
rect 33140 6196 33192 6248
rect 34796 6196 34848 6248
rect 36084 6196 36136 6248
rect 37924 6196 37976 6248
rect 39856 6273 39865 6307
rect 39865 6273 39899 6307
rect 39899 6273 39908 6307
rect 39856 6264 39908 6273
rect 40408 6307 40460 6316
rect 40408 6273 40417 6307
rect 40417 6273 40451 6307
rect 40451 6273 40460 6307
rect 40408 6264 40460 6273
rect 40960 6400 41012 6452
rect 41512 6400 41564 6452
rect 43904 6443 43956 6452
rect 43904 6409 43913 6443
rect 43913 6409 43947 6443
rect 43947 6409 43956 6443
rect 43904 6400 43956 6409
rect 45008 6400 45060 6452
rect 49884 6443 49936 6452
rect 49884 6409 49893 6443
rect 49893 6409 49927 6443
rect 49927 6409 49936 6443
rect 49884 6400 49936 6409
rect 50344 6400 50396 6452
rect 51540 6400 51592 6452
rect 46848 6332 46900 6384
rect 47584 6332 47636 6384
rect 49148 6332 49200 6384
rect 41052 6264 41104 6316
rect 42524 6264 42576 6316
rect 41144 6196 41196 6248
rect 46296 6307 46348 6316
rect 44916 6196 44968 6248
rect 28816 6128 28868 6180
rect 35440 6128 35492 6180
rect 38660 6128 38712 6180
rect 38844 6128 38896 6180
rect 25044 6060 25096 6112
rect 27896 6103 27948 6112
rect 27896 6069 27905 6103
rect 27905 6069 27939 6103
rect 27939 6069 27948 6103
rect 27896 6060 27948 6069
rect 27988 6060 28040 6112
rect 28448 6060 28500 6112
rect 33968 6060 34020 6112
rect 36176 6060 36228 6112
rect 36636 6060 36688 6112
rect 38016 6060 38068 6112
rect 38292 6060 38344 6112
rect 39856 6060 39908 6112
rect 42616 6060 42668 6112
rect 44640 6060 44692 6112
rect 46296 6273 46305 6307
rect 46305 6273 46339 6307
rect 46339 6273 46348 6307
rect 46296 6264 46348 6273
rect 46388 6264 46440 6316
rect 46756 6307 46808 6316
rect 46756 6273 46765 6307
rect 46765 6273 46799 6307
rect 46799 6273 46808 6307
rect 46756 6264 46808 6273
rect 47032 6264 47084 6316
rect 48044 6307 48096 6316
rect 48044 6273 48053 6307
rect 48053 6273 48087 6307
rect 48087 6273 48096 6307
rect 48044 6264 48096 6273
rect 48596 6264 48648 6316
rect 50804 6332 50856 6384
rect 51448 6332 51500 6384
rect 49884 6196 49936 6248
rect 47308 6128 47360 6180
rect 45928 6060 45980 6112
rect 49792 6060 49844 6112
rect 50160 6307 50212 6316
rect 50160 6273 50169 6307
rect 50169 6273 50203 6307
rect 50203 6273 50212 6307
rect 50344 6307 50396 6316
rect 50160 6264 50212 6273
rect 50344 6273 50353 6307
rect 50353 6273 50387 6307
rect 50387 6273 50396 6307
rect 50344 6264 50396 6273
rect 50712 6264 50764 6316
rect 51172 6307 51224 6316
rect 51172 6273 51181 6307
rect 51181 6273 51215 6307
rect 51215 6273 51224 6307
rect 51172 6264 51224 6273
rect 53288 6400 53340 6452
rect 54852 6400 54904 6452
rect 58440 6400 58492 6452
rect 52184 6375 52236 6384
rect 52184 6341 52193 6375
rect 52193 6341 52227 6375
rect 52227 6341 52236 6375
rect 52184 6332 52236 6341
rect 52276 6332 52328 6384
rect 52736 6332 52788 6384
rect 50436 6196 50488 6248
rect 50068 6128 50120 6180
rect 51724 6264 51776 6316
rect 53104 6307 53156 6316
rect 53104 6273 53113 6307
rect 53113 6273 53147 6307
rect 53147 6273 53156 6307
rect 53104 6264 53156 6273
rect 55128 6332 55180 6384
rect 57520 6375 57572 6384
rect 57520 6341 57529 6375
rect 57529 6341 57563 6375
rect 57563 6341 57572 6375
rect 57520 6332 57572 6341
rect 58348 6332 58400 6384
rect 52184 6196 52236 6248
rect 52460 6196 52512 6248
rect 52920 6239 52972 6248
rect 52920 6205 52929 6239
rect 52929 6205 52963 6239
rect 52963 6205 52972 6239
rect 52920 6196 52972 6205
rect 53012 6196 53064 6248
rect 54208 6196 54260 6248
rect 51540 6128 51592 6180
rect 53840 6128 53892 6180
rect 56508 6128 56560 6180
rect 53472 6060 53524 6112
rect 54116 6060 54168 6112
rect 56600 6060 56652 6112
rect 56876 6103 56928 6112
rect 56876 6069 56885 6103
rect 56885 6069 56919 6103
rect 56919 6069 56928 6103
rect 56876 6060 56928 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2412 5899 2464 5908
rect 2412 5865 2421 5899
rect 2421 5865 2455 5899
rect 2455 5865 2464 5899
rect 2412 5856 2464 5865
rect 25872 5899 25924 5908
rect 25872 5865 25881 5899
rect 25881 5865 25915 5899
rect 25915 5865 25924 5899
rect 25872 5856 25924 5865
rect 27160 5899 27212 5908
rect 27160 5865 27169 5899
rect 27169 5865 27203 5899
rect 27203 5865 27212 5899
rect 27160 5856 27212 5865
rect 25780 5788 25832 5840
rect 28724 5856 28776 5908
rect 31392 5899 31444 5908
rect 31392 5865 31401 5899
rect 31401 5865 31435 5899
rect 31435 5865 31444 5899
rect 31392 5856 31444 5865
rect 27620 5720 27672 5772
rect 2412 5652 2464 5704
rect 26056 5695 26108 5704
rect 26056 5661 26065 5695
rect 26065 5661 26099 5695
rect 26099 5661 26108 5695
rect 26056 5652 26108 5661
rect 27344 5695 27396 5704
rect 26424 5627 26476 5636
rect 26424 5593 26433 5627
rect 26433 5593 26467 5627
rect 26467 5593 26476 5627
rect 26424 5584 26476 5593
rect 27344 5661 27350 5695
rect 27350 5661 27384 5695
rect 27384 5661 27396 5695
rect 27344 5652 27396 5661
rect 27712 5695 27764 5704
rect 27712 5661 27721 5695
rect 27721 5661 27755 5695
rect 27755 5661 27764 5695
rect 27712 5652 27764 5661
rect 28632 5788 28684 5840
rect 29552 5788 29604 5840
rect 30748 5788 30800 5840
rect 32220 5856 32272 5908
rect 34060 5899 34112 5908
rect 32956 5788 33008 5840
rect 32036 5720 32088 5772
rect 32588 5763 32640 5772
rect 32588 5729 32597 5763
rect 32597 5729 32631 5763
rect 32631 5729 32640 5763
rect 32588 5720 32640 5729
rect 33140 5763 33192 5772
rect 33140 5729 33149 5763
rect 33149 5729 33183 5763
rect 33183 5729 33192 5763
rect 33140 5720 33192 5729
rect 34060 5865 34069 5899
rect 34069 5865 34103 5899
rect 34103 5865 34112 5899
rect 34060 5856 34112 5865
rect 34428 5856 34480 5908
rect 35624 5856 35676 5908
rect 28632 5652 28684 5704
rect 29644 5652 29696 5704
rect 28540 5584 28592 5636
rect 30196 5695 30248 5704
rect 30196 5661 30205 5695
rect 30205 5661 30239 5695
rect 30239 5661 30248 5695
rect 30196 5652 30248 5661
rect 30564 5652 30616 5704
rect 31852 5695 31904 5704
rect 31852 5661 31861 5695
rect 31861 5661 31895 5695
rect 31895 5661 31904 5695
rect 31852 5652 31904 5661
rect 33048 5584 33100 5636
rect 33232 5584 33284 5636
rect 35164 5720 35216 5772
rect 34244 5652 34296 5704
rect 35348 5720 35400 5772
rect 36912 5788 36964 5840
rect 39488 5856 39540 5908
rect 42156 5899 42208 5908
rect 42156 5865 42165 5899
rect 42165 5865 42199 5899
rect 42199 5865 42208 5899
rect 42156 5856 42208 5865
rect 42800 5856 42852 5908
rect 46204 5856 46256 5908
rect 40684 5788 40736 5840
rect 41420 5788 41472 5840
rect 36360 5763 36412 5772
rect 36360 5729 36369 5763
rect 36369 5729 36403 5763
rect 36403 5729 36412 5763
rect 37004 5763 37056 5772
rect 36360 5720 36412 5729
rect 37004 5729 37013 5763
rect 37013 5729 37047 5763
rect 37047 5729 37056 5763
rect 37004 5720 37056 5729
rect 36176 5652 36228 5704
rect 38016 5695 38068 5704
rect 38016 5661 38025 5695
rect 38025 5661 38059 5695
rect 38059 5661 38068 5695
rect 38016 5652 38068 5661
rect 38200 5695 38252 5704
rect 38200 5661 38217 5695
rect 38217 5661 38252 5695
rect 38200 5652 38252 5661
rect 38292 5695 38344 5704
rect 38292 5661 38301 5695
rect 38301 5661 38335 5695
rect 38335 5661 38344 5695
rect 38292 5652 38344 5661
rect 38476 5695 38528 5704
rect 38476 5661 38485 5695
rect 38485 5661 38519 5695
rect 38519 5661 38528 5695
rect 38476 5652 38528 5661
rect 39120 5652 39172 5704
rect 39396 5652 39448 5704
rect 40040 5652 40092 5704
rect 41144 5652 41196 5704
rect 41328 5695 41380 5704
rect 41328 5661 41337 5695
rect 41337 5661 41371 5695
rect 41371 5661 41380 5695
rect 41328 5652 41380 5661
rect 34612 5584 34664 5636
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 27344 5559 27396 5568
rect 27344 5525 27353 5559
rect 27353 5525 27387 5559
rect 27387 5525 27396 5559
rect 27344 5516 27396 5525
rect 28356 5516 28408 5568
rect 28724 5516 28776 5568
rect 29552 5516 29604 5568
rect 34704 5516 34756 5568
rect 35072 5559 35124 5568
rect 35072 5525 35081 5559
rect 35081 5525 35115 5559
rect 35115 5525 35124 5559
rect 35072 5516 35124 5525
rect 35256 5516 35308 5568
rect 37004 5584 37056 5636
rect 35716 5516 35768 5568
rect 41236 5584 41288 5636
rect 43168 5720 43220 5772
rect 43352 5763 43404 5772
rect 43352 5729 43361 5763
rect 43361 5729 43395 5763
rect 43395 5729 43404 5763
rect 43352 5720 43404 5729
rect 45284 5763 45336 5772
rect 45284 5729 45293 5763
rect 45293 5729 45327 5763
rect 45327 5729 45336 5763
rect 45284 5720 45336 5729
rect 46388 5720 46440 5772
rect 48780 5856 48832 5908
rect 50436 5856 50488 5908
rect 50988 5856 51040 5908
rect 48320 5831 48372 5840
rect 48320 5797 48329 5831
rect 48329 5797 48363 5831
rect 48363 5797 48372 5831
rect 48320 5788 48372 5797
rect 50620 5831 50672 5840
rect 50620 5797 50629 5831
rect 50629 5797 50663 5831
rect 50663 5797 50672 5831
rect 50620 5788 50672 5797
rect 52368 5856 52420 5908
rect 52920 5856 52972 5908
rect 53564 5856 53616 5908
rect 56508 5856 56560 5908
rect 57152 5899 57204 5908
rect 57152 5865 57161 5899
rect 57161 5865 57195 5899
rect 57195 5865 57204 5899
rect 57152 5856 57204 5865
rect 58532 5856 58584 5908
rect 55496 5831 55548 5840
rect 43260 5695 43312 5704
rect 43260 5661 43269 5695
rect 43269 5661 43303 5695
rect 43303 5661 43312 5695
rect 43260 5652 43312 5661
rect 42064 5584 42116 5636
rect 42984 5584 43036 5636
rect 44272 5627 44324 5636
rect 44272 5593 44281 5627
rect 44281 5593 44315 5627
rect 44315 5593 44324 5627
rect 44272 5584 44324 5593
rect 44916 5584 44968 5636
rect 45468 5652 45520 5704
rect 40684 5516 40736 5568
rect 41052 5559 41104 5568
rect 41052 5525 41061 5559
rect 41061 5525 41095 5559
rect 41095 5525 41104 5559
rect 41052 5516 41104 5525
rect 42340 5516 42392 5568
rect 43996 5516 44048 5568
rect 45652 5627 45704 5636
rect 45652 5593 45661 5627
rect 45661 5593 45695 5627
rect 45695 5593 45704 5627
rect 47216 5652 47268 5704
rect 47768 5652 47820 5704
rect 48044 5695 48096 5704
rect 48044 5661 48053 5695
rect 48053 5661 48087 5695
rect 48087 5661 48096 5695
rect 48044 5652 48096 5661
rect 45652 5584 45704 5593
rect 47492 5584 47544 5636
rect 48780 5720 48832 5772
rect 49884 5720 49936 5772
rect 55496 5797 55505 5831
rect 55505 5797 55539 5831
rect 55539 5797 55548 5831
rect 55496 5788 55548 5797
rect 51908 5720 51960 5772
rect 53104 5763 53156 5772
rect 53104 5729 53113 5763
rect 53113 5729 53147 5763
rect 53147 5729 53156 5763
rect 53104 5720 53156 5729
rect 54116 5763 54168 5772
rect 54116 5729 54125 5763
rect 54125 5729 54159 5763
rect 54159 5729 54168 5763
rect 54116 5720 54168 5729
rect 54760 5720 54812 5772
rect 55036 5720 55088 5772
rect 48596 5695 48648 5704
rect 48596 5661 48605 5695
rect 48605 5661 48639 5695
rect 48639 5661 48648 5695
rect 48596 5652 48648 5661
rect 49608 5652 49660 5704
rect 50896 5652 50948 5704
rect 48688 5584 48740 5636
rect 53472 5652 53524 5704
rect 54208 5695 54260 5704
rect 54208 5661 54217 5695
rect 54217 5661 54251 5695
rect 54251 5661 54260 5695
rect 54208 5652 54260 5661
rect 54852 5695 54904 5704
rect 54852 5661 54861 5695
rect 54861 5661 54895 5695
rect 54895 5661 54904 5695
rect 54852 5652 54904 5661
rect 55128 5584 55180 5636
rect 45744 5516 45796 5568
rect 46020 5516 46072 5568
rect 46940 5516 46992 5568
rect 52920 5516 52972 5568
rect 54852 5559 54904 5568
rect 54852 5525 54861 5559
rect 54861 5525 54895 5559
rect 54895 5525 54904 5559
rect 54852 5516 54904 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 26148 5355 26200 5364
rect 26148 5321 26157 5355
rect 26157 5321 26191 5355
rect 26191 5321 26200 5355
rect 26148 5312 26200 5321
rect 27344 5355 27396 5364
rect 27344 5321 27353 5355
rect 27353 5321 27387 5355
rect 27387 5321 27396 5355
rect 27344 5312 27396 5321
rect 25964 5244 26016 5296
rect 28816 5312 28868 5364
rect 30104 5355 30156 5364
rect 30104 5321 30113 5355
rect 30113 5321 30147 5355
rect 30147 5321 30156 5355
rect 30104 5312 30156 5321
rect 31852 5312 31904 5364
rect 33048 5312 33100 5364
rect 33784 5355 33836 5364
rect 33784 5321 33793 5355
rect 33793 5321 33827 5355
rect 33827 5321 33836 5355
rect 33784 5312 33836 5321
rect 26332 5176 26384 5228
rect 26792 5176 26844 5228
rect 27804 5219 27856 5228
rect 26976 5108 27028 5160
rect 27804 5185 27813 5219
rect 27813 5185 27847 5219
rect 27847 5185 27856 5219
rect 27804 5176 27856 5185
rect 29368 5176 29420 5228
rect 29552 5219 29604 5228
rect 29552 5185 29561 5219
rect 29561 5185 29595 5219
rect 29595 5185 29604 5219
rect 29552 5176 29604 5185
rect 30196 5244 30248 5296
rect 29184 5108 29236 5160
rect 30748 5176 30800 5228
rect 31300 5219 31352 5228
rect 31300 5185 31309 5219
rect 31309 5185 31343 5219
rect 31343 5185 31352 5219
rect 31300 5176 31352 5185
rect 32312 5244 32364 5296
rect 32496 5244 32548 5296
rect 35808 5244 35860 5296
rect 31484 5219 31536 5228
rect 31484 5185 31493 5219
rect 31493 5185 31527 5219
rect 31527 5185 31536 5219
rect 31484 5176 31536 5185
rect 31852 5176 31904 5228
rect 32680 5176 32732 5228
rect 37648 5244 37700 5296
rect 38200 5244 38252 5296
rect 40040 5244 40092 5296
rect 41052 5244 41104 5296
rect 41788 5244 41840 5296
rect 42800 5244 42852 5296
rect 27988 5040 28040 5092
rect 28264 5040 28316 5092
rect 30472 5040 30524 5092
rect 33232 5151 33284 5160
rect 33232 5117 33241 5151
rect 33241 5117 33275 5151
rect 33275 5117 33284 5151
rect 33232 5108 33284 5117
rect 33416 5108 33468 5160
rect 34520 5151 34572 5160
rect 34520 5117 34529 5151
rect 34529 5117 34563 5151
rect 34563 5117 34572 5151
rect 34520 5108 34572 5117
rect 37188 5108 37240 5160
rect 32772 5040 32824 5092
rect 26884 4972 26936 5024
rect 28908 5015 28960 5024
rect 28908 4981 28917 5015
rect 28917 4981 28951 5015
rect 28951 4981 28960 5015
rect 28908 4972 28960 4981
rect 30196 4972 30248 5024
rect 32312 4972 32364 5024
rect 37924 5219 37976 5228
rect 37924 5185 37933 5219
rect 37933 5185 37967 5219
rect 37967 5185 37976 5219
rect 37924 5176 37976 5185
rect 38476 5176 38528 5228
rect 41420 5176 41472 5228
rect 46664 5312 46716 5364
rect 46848 5355 46900 5364
rect 46848 5321 46857 5355
rect 46857 5321 46891 5355
rect 46891 5321 46900 5355
rect 46848 5312 46900 5321
rect 47492 5312 47544 5364
rect 49700 5312 49752 5364
rect 50804 5312 50856 5364
rect 54116 5312 54168 5364
rect 54852 5312 54904 5364
rect 55312 5312 55364 5364
rect 43720 5244 43772 5296
rect 45560 5244 45612 5296
rect 47860 5287 47912 5296
rect 44640 5219 44692 5228
rect 44640 5185 44649 5219
rect 44649 5185 44683 5219
rect 44683 5185 44692 5219
rect 44640 5176 44692 5185
rect 45284 5176 45336 5228
rect 47032 5219 47084 5228
rect 47032 5185 47041 5219
rect 47041 5185 47075 5219
rect 47075 5185 47084 5219
rect 47032 5176 47084 5185
rect 47860 5253 47869 5287
rect 47869 5253 47903 5287
rect 47903 5253 47912 5287
rect 47860 5244 47912 5253
rect 50528 5244 50580 5296
rect 53748 5244 53800 5296
rect 55128 5244 55180 5296
rect 57980 5244 58032 5296
rect 48596 5176 48648 5228
rect 49332 5219 49384 5228
rect 38016 5108 38068 5160
rect 38568 5151 38620 5160
rect 38568 5117 38577 5151
rect 38577 5117 38611 5151
rect 38611 5117 38620 5151
rect 38568 5108 38620 5117
rect 40592 5151 40644 5160
rect 40592 5117 40601 5151
rect 40601 5117 40635 5151
rect 40635 5117 40644 5151
rect 40592 5108 40644 5117
rect 40960 5108 41012 5160
rect 41604 5108 41656 5160
rect 42064 5108 42116 5160
rect 38936 5040 38988 5092
rect 40776 5040 40828 5092
rect 45836 5108 45888 5160
rect 49056 5108 49108 5160
rect 48504 5040 48556 5092
rect 49332 5185 49341 5219
rect 49341 5185 49375 5219
rect 49375 5185 49384 5219
rect 49332 5176 49384 5185
rect 51632 5219 51684 5228
rect 51632 5185 51641 5219
rect 51641 5185 51675 5219
rect 51675 5185 51684 5219
rect 51632 5176 51684 5185
rect 52276 5176 52328 5228
rect 53472 5176 53524 5228
rect 49240 5108 49292 5160
rect 49608 5108 49660 5160
rect 56048 5176 56100 5228
rect 54668 5108 54720 5160
rect 57520 5108 57572 5160
rect 37280 4972 37332 5024
rect 40500 4972 40552 5024
rect 41604 4972 41656 5024
rect 46204 4972 46256 5024
rect 46480 4972 46532 5024
rect 48596 4972 48648 5024
rect 48780 5015 48832 5024
rect 48780 4981 48789 5015
rect 48789 4981 48823 5015
rect 48823 4981 48832 5015
rect 48780 4972 48832 4981
rect 50620 5040 50672 5092
rect 50804 5015 50856 5024
rect 50804 4981 50813 5015
rect 50813 4981 50847 5015
rect 50847 4981 50856 5015
rect 50804 4972 50856 4981
rect 51632 4972 51684 5024
rect 55036 4972 55088 5024
rect 56508 5015 56560 5024
rect 56508 4981 56517 5015
rect 56517 4981 56551 5015
rect 56551 4981 56560 5015
rect 56508 4972 56560 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 26056 4768 26108 4820
rect 27252 4811 27304 4820
rect 27252 4777 27261 4811
rect 27261 4777 27295 4811
rect 27295 4777 27304 4811
rect 27252 4768 27304 4777
rect 27712 4768 27764 4820
rect 29368 4768 29420 4820
rect 30012 4768 30064 4820
rect 31116 4768 31168 4820
rect 32496 4811 32548 4820
rect 32496 4777 32505 4811
rect 32505 4777 32539 4811
rect 32539 4777 32548 4811
rect 32496 4768 32548 4777
rect 33048 4768 33100 4820
rect 33692 4768 33744 4820
rect 34152 4768 34204 4820
rect 37556 4768 37608 4820
rect 37832 4768 37884 4820
rect 41328 4768 41380 4820
rect 41880 4768 41932 4820
rect 42432 4768 42484 4820
rect 45744 4768 45796 4820
rect 45836 4811 45888 4820
rect 45836 4777 45845 4811
rect 45845 4777 45879 4811
rect 45879 4777 45888 4811
rect 45836 4768 45888 4777
rect 47400 4811 47452 4820
rect 47400 4777 47409 4811
rect 47409 4777 47443 4811
rect 47443 4777 47452 4811
rect 47400 4768 47452 4777
rect 47676 4768 47728 4820
rect 51540 4811 51592 4820
rect 51540 4777 51549 4811
rect 51549 4777 51583 4811
rect 51583 4777 51592 4811
rect 51540 4768 51592 4777
rect 52828 4768 52880 4820
rect 54024 4768 54076 4820
rect 56048 4811 56100 4820
rect 56048 4777 56057 4811
rect 56057 4777 56091 4811
rect 56091 4777 56100 4811
rect 56048 4768 56100 4777
rect 26332 4700 26384 4752
rect 28816 4700 28868 4752
rect 27804 4632 27856 4684
rect 28356 4632 28408 4684
rect 31208 4700 31260 4752
rect 31852 4743 31904 4752
rect 31852 4709 31861 4743
rect 31861 4709 31895 4743
rect 31895 4709 31904 4743
rect 31852 4700 31904 4709
rect 30196 4675 30248 4684
rect 30196 4641 30205 4675
rect 30205 4641 30239 4675
rect 30239 4641 30248 4675
rect 30196 4632 30248 4641
rect 34612 4700 34664 4752
rect 38568 4700 38620 4752
rect 42524 4700 42576 4752
rect 43628 4700 43680 4752
rect 47768 4700 47820 4752
rect 33416 4632 33468 4684
rect 33784 4632 33836 4684
rect 33876 4632 33928 4684
rect 37096 4632 37148 4684
rect 37464 4632 37516 4684
rect 28080 4564 28132 4616
rect 28264 4607 28316 4616
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 28448 4607 28500 4616
rect 28448 4573 28457 4607
rect 28457 4573 28491 4607
rect 28491 4573 28500 4607
rect 28448 4564 28500 4573
rect 25320 4496 25372 4548
rect 29092 4564 29144 4616
rect 29828 4564 29880 4616
rect 31484 4564 31536 4616
rect 32312 4564 32364 4616
rect 32864 4607 32916 4616
rect 32864 4573 32873 4607
rect 32873 4573 32907 4607
rect 32907 4573 32916 4607
rect 32864 4564 32916 4573
rect 38108 4564 38160 4616
rect 40224 4632 40276 4684
rect 41696 4632 41748 4684
rect 41880 4564 41932 4616
rect 42156 4632 42208 4684
rect 42432 4632 42484 4684
rect 45192 4675 45244 4684
rect 45192 4641 45201 4675
rect 45201 4641 45235 4675
rect 45235 4641 45244 4675
rect 45192 4632 45244 4641
rect 45744 4632 45796 4684
rect 48872 4632 48924 4684
rect 49332 4632 49384 4684
rect 42064 4564 42116 4616
rect 31208 4496 31260 4548
rect 28172 4428 28224 4480
rect 35348 4539 35400 4548
rect 33876 4428 33928 4480
rect 34060 4428 34112 4480
rect 35348 4505 35357 4539
rect 35357 4505 35391 4539
rect 35391 4505 35400 4539
rect 35348 4496 35400 4505
rect 36084 4496 36136 4548
rect 37096 4496 37148 4548
rect 42340 4496 42392 4548
rect 37648 4428 37700 4480
rect 40684 4471 40736 4480
rect 40684 4437 40693 4471
rect 40693 4437 40727 4471
rect 40727 4437 40736 4471
rect 40684 4428 40736 4437
rect 41512 4428 41564 4480
rect 42892 4607 42944 4616
rect 42892 4573 42901 4607
rect 42901 4573 42935 4607
rect 42935 4573 42944 4607
rect 46940 4607 46992 4616
rect 42892 4564 42944 4573
rect 43444 4539 43496 4548
rect 43444 4505 43453 4539
rect 43453 4505 43487 4539
rect 43487 4505 43496 4539
rect 43444 4496 43496 4505
rect 43536 4496 43588 4548
rect 45192 4496 45244 4548
rect 46020 4496 46072 4548
rect 44180 4428 44232 4480
rect 45652 4428 45704 4480
rect 45928 4428 45980 4480
rect 46388 4428 46440 4480
rect 46940 4573 46949 4607
rect 46949 4573 46983 4607
rect 46983 4573 46992 4607
rect 49976 4700 50028 4752
rect 50804 4632 50856 4684
rect 53104 4700 53156 4752
rect 55220 4700 55272 4752
rect 54208 4632 54260 4684
rect 46940 4564 46992 4573
rect 50160 4564 50212 4616
rect 50528 4564 50580 4616
rect 54576 4564 54628 4616
rect 55588 4564 55640 4616
rect 46664 4496 46716 4548
rect 48044 4496 48096 4548
rect 52000 4496 52052 4548
rect 47308 4428 47360 4480
rect 47492 4428 47544 4480
rect 48596 4428 48648 4480
rect 49608 4471 49660 4480
rect 49608 4437 49617 4471
rect 49617 4437 49651 4471
rect 49651 4437 49660 4471
rect 49608 4428 49660 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 28448 4224 28500 4276
rect 31852 4224 31904 4276
rect 32772 4224 32824 4276
rect 33876 4224 33928 4276
rect 34060 4267 34112 4276
rect 34060 4233 34069 4267
rect 34069 4233 34103 4267
rect 34103 4233 34112 4267
rect 34060 4224 34112 4233
rect 34152 4267 34204 4276
rect 34152 4233 34161 4267
rect 34161 4233 34195 4267
rect 34195 4233 34204 4267
rect 34152 4224 34204 4233
rect 34796 4224 34848 4276
rect 35808 4224 35860 4276
rect 29092 4199 29144 4208
rect 29092 4165 29101 4199
rect 29101 4165 29135 4199
rect 29135 4165 29144 4199
rect 29092 4156 29144 4165
rect 29828 4156 29880 4208
rect 32404 4199 32456 4208
rect 32404 4165 32413 4199
rect 32413 4165 32447 4199
rect 32447 4165 32456 4199
rect 32404 4156 32456 4165
rect 28080 4088 28132 4140
rect 28356 4131 28408 4140
rect 28356 4097 28365 4131
rect 28365 4097 28399 4131
rect 28399 4097 28408 4131
rect 28356 4088 28408 4097
rect 30196 4131 30248 4140
rect 27988 4063 28040 4072
rect 27988 4029 27997 4063
rect 27997 4029 28031 4063
rect 28031 4029 28040 4063
rect 27988 4020 28040 4029
rect 30196 4097 30205 4131
rect 30205 4097 30239 4131
rect 30239 4097 30248 4131
rect 30196 4088 30248 4097
rect 30288 4088 30340 4140
rect 31484 4088 31536 4140
rect 32220 4020 32272 4072
rect 32496 4131 32548 4140
rect 32496 4097 32505 4131
rect 32505 4097 32539 4131
rect 32539 4097 32548 4131
rect 32496 4088 32548 4097
rect 32680 4131 32732 4140
rect 32680 4097 32689 4131
rect 32689 4097 32723 4131
rect 32723 4097 32732 4131
rect 32680 4088 32732 4097
rect 33968 4088 34020 4140
rect 32588 4020 32640 4072
rect 34152 4020 34204 4072
rect 34704 4156 34756 4208
rect 37096 4224 37148 4276
rect 37280 4156 37332 4208
rect 40868 4224 40920 4276
rect 43628 4224 43680 4276
rect 46204 4224 46256 4276
rect 40040 4156 40092 4208
rect 40316 4156 40368 4208
rect 41696 4156 41748 4208
rect 43536 4156 43588 4208
rect 43720 4156 43772 4208
rect 45008 4199 45060 4208
rect 45008 4165 45010 4199
rect 45010 4165 45044 4199
rect 45044 4165 45060 4199
rect 45008 4156 45060 4165
rect 47584 4156 47636 4208
rect 41144 4088 41196 4140
rect 42616 4131 42668 4140
rect 42616 4097 42625 4131
rect 42625 4097 42659 4131
rect 42659 4097 42668 4131
rect 42616 4088 42668 4097
rect 43352 4088 43404 4140
rect 45284 4131 45336 4140
rect 45284 4097 45293 4131
rect 45293 4097 45327 4131
rect 45327 4097 45336 4131
rect 45744 4131 45796 4140
rect 45284 4088 45336 4097
rect 45744 4097 45753 4131
rect 45753 4097 45787 4131
rect 45787 4097 45796 4131
rect 45744 4088 45796 4097
rect 48964 4199 49016 4208
rect 48964 4165 48973 4199
rect 48973 4165 49007 4199
rect 49007 4165 49016 4199
rect 48964 4156 49016 4165
rect 49608 4156 49660 4208
rect 52552 4156 52604 4208
rect 53104 4199 53156 4208
rect 53104 4165 53113 4199
rect 53113 4165 53147 4199
rect 53147 4165 53156 4199
rect 53104 4156 53156 4165
rect 54208 4224 54260 4276
rect 55128 4224 55180 4276
rect 54944 4156 54996 4208
rect 55496 4156 55548 4208
rect 27804 3952 27856 4004
rect 29460 3952 29512 4004
rect 30288 3884 30340 3936
rect 33876 3952 33928 4004
rect 31852 3884 31904 3936
rect 33048 3884 33100 3936
rect 37280 4020 37332 4072
rect 37464 4063 37516 4072
rect 37464 4029 37473 4063
rect 37473 4029 37507 4063
rect 37507 4029 37516 4063
rect 37464 4020 37516 4029
rect 37740 4063 37792 4072
rect 37740 4029 37749 4063
rect 37749 4029 37783 4063
rect 37783 4029 37792 4063
rect 37740 4020 37792 4029
rect 38476 4020 38528 4072
rect 40040 4063 40092 4072
rect 40040 4029 40049 4063
rect 40049 4029 40083 4063
rect 40083 4029 40092 4063
rect 40040 4020 40092 4029
rect 41512 3995 41564 4004
rect 37372 3884 37424 3936
rect 41512 3961 41521 3995
rect 41521 3961 41555 3995
rect 41555 3961 41564 3995
rect 41512 3952 41564 3961
rect 45560 3952 45612 4004
rect 48136 3952 48188 4004
rect 49884 4088 49936 4140
rect 50896 4088 50948 4140
rect 54208 4020 54260 4072
rect 50712 3952 50764 4004
rect 52184 3952 52236 4004
rect 54668 3952 54720 4004
rect 38292 3884 38344 3936
rect 43352 3884 43404 3936
rect 43444 3884 43496 3936
rect 45652 3884 45704 3936
rect 46480 3884 46532 3936
rect 48228 3884 48280 3936
rect 51172 3927 51224 3936
rect 51172 3893 51181 3927
rect 51181 3893 51215 3927
rect 51215 3893 51224 3927
rect 51172 3884 51224 3893
rect 53472 3884 53524 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 28448 3680 28500 3732
rect 29736 3723 29788 3732
rect 29736 3689 29745 3723
rect 29745 3689 29779 3723
rect 29779 3689 29788 3723
rect 29736 3680 29788 3689
rect 30012 3680 30064 3732
rect 31300 3723 31352 3732
rect 31300 3689 31309 3723
rect 31309 3689 31343 3723
rect 31343 3689 31352 3723
rect 31300 3680 31352 3689
rect 31852 3723 31904 3732
rect 31852 3689 31861 3723
rect 31861 3689 31895 3723
rect 31895 3689 31904 3723
rect 31852 3680 31904 3689
rect 32220 3680 32272 3732
rect 33692 3680 33744 3732
rect 37188 3680 37240 3732
rect 32680 3612 32732 3664
rect 32864 3612 32916 3664
rect 34060 3612 34112 3664
rect 36268 3612 36320 3664
rect 40040 3680 40092 3732
rect 43352 3680 43404 3732
rect 47584 3723 47636 3732
rect 45744 3612 45796 3664
rect 30288 3544 30340 3596
rect 30196 3476 30248 3528
rect 32496 3476 32548 3528
rect 32588 3519 32640 3528
rect 32588 3485 32609 3519
rect 32609 3485 32640 3519
rect 33968 3544 34020 3596
rect 34336 3544 34388 3596
rect 32588 3476 32640 3485
rect 33876 3476 33928 3528
rect 34060 3476 34112 3528
rect 31208 3340 31260 3392
rect 33600 3408 33652 3460
rect 34244 3408 34296 3460
rect 37280 3544 37332 3596
rect 40592 3544 40644 3596
rect 41236 3587 41288 3596
rect 41236 3553 41245 3587
rect 41245 3553 41279 3587
rect 41279 3553 41288 3587
rect 41236 3544 41288 3553
rect 42616 3544 42668 3596
rect 45284 3544 45336 3596
rect 46480 3544 46532 3596
rect 40316 3476 40368 3528
rect 40500 3519 40552 3528
rect 40500 3485 40509 3519
rect 40509 3485 40543 3519
rect 40543 3485 40552 3519
rect 40500 3476 40552 3485
rect 43536 3519 43588 3528
rect 43536 3485 43545 3519
rect 43545 3485 43579 3519
rect 43579 3485 43588 3519
rect 43536 3476 43588 3485
rect 43812 3476 43864 3528
rect 34612 3340 34664 3392
rect 35716 3408 35768 3460
rect 37096 3408 37148 3460
rect 36360 3340 36412 3392
rect 37464 3408 37516 3460
rect 43720 3451 43772 3460
rect 43720 3417 43729 3451
rect 43729 3417 43763 3451
rect 43763 3417 43772 3451
rect 43720 3408 43772 3417
rect 46664 3408 46716 3460
rect 47584 3689 47593 3723
rect 47593 3689 47627 3723
rect 47627 3689 47636 3723
rect 47584 3680 47636 3689
rect 50068 3680 50120 3732
rect 54208 3680 54260 3732
rect 54668 3723 54720 3732
rect 54668 3689 54677 3723
rect 54677 3689 54711 3723
rect 54711 3689 54720 3723
rect 54668 3680 54720 3689
rect 55496 3723 55548 3732
rect 55496 3689 55505 3723
rect 55505 3689 55539 3723
rect 55539 3689 55548 3723
rect 55496 3680 55548 3689
rect 47860 3612 47912 3664
rect 49240 3655 49292 3664
rect 49240 3621 49249 3655
rect 49249 3621 49283 3655
rect 49283 3621 49292 3655
rect 49240 3612 49292 3621
rect 51172 3612 51224 3664
rect 56508 3612 56560 3664
rect 48872 3519 48924 3528
rect 48872 3485 48881 3519
rect 48881 3485 48915 3519
rect 48915 3485 48924 3519
rect 48872 3476 48924 3485
rect 51448 3476 51500 3528
rect 51356 3408 51408 3460
rect 52000 3408 52052 3460
rect 40132 3340 40184 3392
rect 44180 3340 44232 3392
rect 45928 3340 45980 3392
rect 49240 3340 49292 3392
rect 52276 3476 52328 3528
rect 53472 3340 53524 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 26424 3136 26476 3188
rect 30196 3111 30248 3120
rect 30196 3077 30205 3111
rect 30205 3077 30239 3111
rect 30239 3077 30248 3111
rect 30196 3068 30248 3077
rect 31208 3068 31260 3120
rect 31484 3111 31536 3120
rect 31484 3077 31493 3111
rect 31493 3077 31527 3111
rect 31527 3077 31536 3111
rect 31484 3068 31536 3077
rect 29184 3043 29236 3052
rect 29184 3009 29193 3043
rect 29193 3009 29227 3043
rect 29227 3009 29236 3043
rect 32680 3068 32732 3120
rect 32864 3068 32916 3120
rect 29184 3000 29236 3009
rect 32036 3000 32088 3052
rect 34336 3136 34388 3188
rect 34520 3136 34572 3188
rect 34796 3068 34848 3120
rect 35440 3068 35492 3120
rect 37280 3136 37332 3188
rect 37648 3136 37700 3188
rect 40316 3136 40368 3188
rect 41788 3179 41840 3188
rect 41788 3145 41797 3179
rect 41797 3145 41831 3179
rect 41831 3145 41840 3179
rect 41788 3136 41840 3145
rect 43720 3136 43772 3188
rect 47768 3179 47820 3188
rect 35716 3068 35768 3120
rect 27896 2932 27948 2984
rect 36268 3000 36320 3052
rect 30472 2864 30524 2916
rect 31208 2907 31260 2916
rect 31208 2873 31217 2907
rect 31217 2873 31251 2907
rect 31251 2873 31260 2907
rect 31208 2864 31260 2873
rect 34244 2864 34296 2916
rect 36452 2864 36504 2916
rect 39304 3068 39356 3120
rect 40408 3068 40460 3120
rect 40592 3068 40644 3120
rect 37280 3000 37332 3052
rect 38476 3000 38528 3052
rect 40868 3000 40920 3052
rect 37556 2932 37608 2984
rect 38108 2932 38160 2984
rect 40224 2932 40276 2984
rect 40776 2975 40828 2984
rect 40776 2941 40785 2975
rect 40785 2941 40819 2975
rect 40819 2941 40828 2975
rect 40776 2932 40828 2941
rect 40960 2932 41012 2984
rect 42984 3068 43036 3120
rect 47768 3145 47777 3179
rect 47777 3145 47811 3179
rect 47811 3145 47820 3179
rect 47768 3136 47820 3145
rect 45284 3068 45336 3120
rect 45376 3111 45428 3120
rect 45376 3077 45385 3111
rect 45385 3077 45419 3111
rect 45419 3077 45428 3111
rect 45376 3068 45428 3077
rect 46664 3068 46716 3120
rect 46756 3068 46808 3120
rect 48136 3068 48188 3120
rect 48412 3111 48464 3120
rect 48412 3077 48421 3111
rect 48421 3077 48455 3111
rect 48455 3077 48464 3111
rect 48412 3068 48464 3077
rect 48780 3068 48832 3120
rect 50896 3136 50948 3188
rect 51448 3136 51500 3188
rect 51908 3136 51960 3188
rect 52276 3136 52328 3188
rect 53472 3179 53524 3188
rect 53472 3145 53481 3179
rect 53481 3145 53515 3179
rect 53515 3145 53524 3179
rect 53472 3136 53524 3145
rect 54208 3136 54260 3188
rect 54576 3179 54628 3188
rect 54576 3145 54585 3179
rect 54585 3145 54619 3179
rect 54619 3145 54628 3179
rect 54576 3136 54628 3145
rect 55220 3179 55272 3188
rect 55220 3145 55229 3179
rect 55229 3145 55263 3179
rect 55263 3145 55272 3179
rect 55220 3136 55272 3145
rect 58164 3136 58216 3188
rect 50160 3111 50212 3120
rect 50160 3077 50169 3111
rect 50169 3077 50203 3111
rect 50203 3077 50212 3111
rect 50160 3068 50212 3077
rect 50712 3111 50764 3120
rect 50712 3077 50721 3111
rect 50721 3077 50755 3111
rect 50755 3077 50764 3111
rect 50712 3068 50764 3077
rect 43260 2932 43312 2984
rect 47216 3000 47268 3052
rect 48228 3000 48280 3052
rect 51356 3000 51408 3052
rect 52184 3000 52236 3052
rect 47124 2975 47176 2984
rect 47124 2941 47133 2975
rect 47133 2941 47167 2975
rect 47167 2941 47176 2975
rect 47124 2932 47176 2941
rect 30288 2796 30340 2848
rect 31024 2796 31076 2848
rect 32312 2796 32364 2848
rect 33692 2796 33744 2848
rect 36360 2796 36412 2848
rect 40040 2796 40092 2848
rect 42892 2796 42944 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 29184 2635 29236 2644
rect 29184 2601 29193 2635
rect 29193 2601 29227 2635
rect 29227 2601 29236 2635
rect 29184 2592 29236 2601
rect 31024 2592 31076 2644
rect 22192 2524 22244 2576
rect 21364 2456 21416 2508
rect 5540 2388 5592 2440
rect 12440 2388 12492 2440
rect 20 2252 72 2304
rect 10968 2252 11020 2304
rect 16764 2252 16816 2304
rect 17684 2295 17736 2304
rect 17684 2261 17693 2295
rect 17693 2261 17727 2295
rect 17727 2261 17736 2295
rect 17684 2252 17736 2261
rect 21916 2252 21968 2304
rect 22836 2295 22888 2304
rect 22836 2261 22845 2295
rect 22845 2261 22879 2295
rect 22879 2261 22888 2295
rect 22836 2252 22888 2261
rect 27712 2252 27764 2304
rect 28908 2388 28960 2440
rect 31300 2592 31352 2644
rect 36268 2592 36320 2644
rect 38108 2592 38160 2644
rect 41328 2592 41380 2644
rect 43168 2592 43220 2644
rect 45192 2592 45244 2644
rect 46204 2592 46256 2644
rect 47032 2635 47084 2644
rect 47032 2601 47041 2635
rect 47041 2601 47075 2635
rect 47075 2601 47084 2635
rect 47032 2592 47084 2601
rect 48688 2592 48740 2644
rect 48872 2635 48924 2644
rect 48872 2601 48881 2635
rect 48881 2601 48915 2635
rect 48915 2601 48924 2635
rect 48872 2592 48924 2601
rect 50896 2592 50948 2644
rect 51632 2635 51684 2644
rect 51632 2601 51641 2635
rect 51641 2601 51675 2635
rect 51675 2601 51684 2635
rect 51632 2592 51684 2601
rect 51908 2592 51960 2644
rect 53472 2635 53524 2644
rect 53472 2601 53481 2635
rect 53481 2601 53515 2635
rect 53515 2601 53524 2635
rect 53472 2592 53524 2601
rect 56968 2635 57020 2644
rect 56968 2601 56977 2635
rect 56977 2601 57011 2635
rect 57011 2601 57020 2635
rect 56968 2592 57020 2601
rect 32496 2524 32548 2576
rect 33876 2524 33928 2576
rect 34796 2524 34848 2576
rect 29920 2388 29972 2440
rect 31208 2431 31260 2440
rect 31208 2397 31217 2431
rect 31217 2397 31251 2431
rect 31251 2397 31260 2431
rect 31208 2388 31260 2397
rect 32680 2388 32732 2440
rect 33140 2388 33192 2440
rect 34152 2431 34204 2440
rect 34152 2397 34161 2431
rect 34161 2397 34195 2431
rect 34195 2397 34204 2431
rect 34152 2388 34204 2397
rect 35348 2388 35400 2440
rect 37464 2499 37516 2508
rect 37464 2465 37473 2499
rect 37473 2465 37507 2499
rect 37507 2465 37516 2499
rect 37464 2456 37516 2465
rect 31300 2252 31352 2304
rect 33508 2320 33560 2372
rect 43536 2524 43588 2576
rect 45652 2524 45704 2576
rect 47124 2524 47176 2576
rect 49240 2524 49292 2576
rect 42248 2456 42300 2508
rect 40040 2431 40092 2440
rect 40040 2397 40049 2431
rect 40049 2397 40083 2431
rect 40083 2397 40092 2431
rect 40040 2388 40092 2397
rect 47032 2388 47084 2440
rect 56968 2388 57020 2440
rect 58164 2388 58216 2440
rect 34428 2252 34480 2304
rect 40684 2320 40736 2372
rect 43536 2320 43588 2372
rect 38660 2252 38712 2304
rect 50160 2252 50212 2304
rect 56048 2252 56100 2304
rect 59912 2252 59964 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 17684 2048 17736 2100
rect 47124 2048 47176 2100
rect 22836 1980 22888 2032
rect 38568 1980 38620 2032
<< metal2 >>
rect 58254 59936 58310 59945
rect 58254 59871 58310 59880
rect 2778 59256 2834 59265
rect 3882 59200 3938 59800
rect 9678 59200 9734 59800
rect 15474 59200 15530 59800
rect 21270 59200 21326 59800
rect 26422 59200 26478 59800
rect 32218 59200 32274 59800
rect 38014 59200 38070 59800
rect 43166 59200 43222 59800
rect 48962 59200 49018 59800
rect 54758 59200 54814 59800
rect 2778 59191 2834 59200
rect 2792 57594 2820 59191
rect 3896 57594 3924 59200
rect 9692 57594 9720 59200
rect 15488 57594 15516 59200
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 21284 57594 21312 59200
rect 26436 57594 26464 59200
rect 2780 57588 2832 57594
rect 2780 57530 2832 57536
rect 3884 57588 3936 57594
rect 3884 57530 3936 57536
rect 9680 57588 9732 57594
rect 9680 57530 9732 57536
rect 15476 57588 15528 57594
rect 15476 57530 15528 57536
rect 21272 57588 21324 57594
rect 21272 57530 21324 57536
rect 26424 57588 26476 57594
rect 26424 57530 26476 57536
rect 28724 57520 28776 57526
rect 28724 57462 28776 57468
rect 2320 57452 2372 57458
rect 2320 57394 2372 57400
rect 4712 57452 4764 57458
rect 4712 57394 4764 57400
rect 10048 57452 10100 57458
rect 10048 57394 10100 57400
rect 15936 57452 15988 57458
rect 15936 57394 15988 57400
rect 22652 57452 22704 57458
rect 22652 57394 22704 57400
rect 27988 57452 28040 57458
rect 27988 57394 28040 57400
rect 2332 57254 2360 57394
rect 4724 57254 4752 57394
rect 2320 57248 2372 57254
rect 2320 57190 2372 57196
rect 4712 57248 4764 57254
rect 4712 57190 4764 57196
rect 1676 53440 1728 53446
rect 1676 53382 1728 53388
rect 1688 53145 1716 53382
rect 1674 53136 1730 53145
rect 1674 53071 1730 53080
rect 1676 47184 1728 47190
rect 1676 47126 1728 47132
rect 1688 47025 1716 47126
rect 1674 47016 1730 47025
rect 1674 46951 1730 46960
rect 1860 41132 1912 41138
rect 1860 41074 1912 41080
rect 1676 40928 1728 40934
rect 1674 40896 1676 40905
rect 1728 40896 1730 40905
rect 1674 40831 1730 40840
rect 1676 35488 1728 35494
rect 1674 35456 1676 35465
rect 1728 35456 1730 35465
rect 1674 35391 1730 35400
rect 1676 29504 1728 29510
rect 1676 29446 1728 29452
rect 1688 29345 1716 29446
rect 1674 29336 1730 29345
rect 1674 29271 1730 29280
rect 1872 29034 1900 41074
rect 1952 35692 2004 35698
rect 1952 35634 2004 35640
rect 1860 29028 1912 29034
rect 1860 28970 1912 28976
rect 1964 25702 1992 35634
rect 1952 25696 2004 25702
rect 1952 25638 2004 25644
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1688 23225 1716 23462
rect 1674 23216 1730 23225
rect 1674 23151 1730 23160
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1596 17814 1624 18226
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1584 17808 1636 17814
rect 1582 17776 1584 17785
rect 1636 17776 1638 17785
rect 1582 17711 1638 17720
rect 1674 11656 1730 11665
rect 1674 11591 1676 11600
rect 1728 11591 1730 11600
rect 1676 11562 1728 11568
rect 1676 5568 1728 5574
rect 1674 5536 1676 5545
rect 1728 5536 1730 5545
rect 1674 5471 1730 5480
rect 1780 5273 1808 18022
rect 1872 12646 1900 23666
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 2332 8294 2360 57190
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 2412 53440 2464 53446
rect 2412 53382 2464 53388
rect 2424 30666 2452 53382
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 2504 46980 2556 46986
rect 2504 46922 2556 46928
rect 2412 30660 2464 30666
rect 2412 30602 2464 30608
rect 2412 29504 2464 29510
rect 2412 29446 2464 29452
rect 2424 27402 2452 29446
rect 2516 28150 2544 46922
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4724 31142 4752 57190
rect 4712 31136 4764 31142
rect 4712 31078 4764 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 2504 28144 2556 28150
rect 2504 28086 2556 28092
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 2412 27396 2464 27402
rect 2412 27338 2464 27344
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 10060 24138 10088 57394
rect 15948 56710 15976 57394
rect 22664 57254 22692 57394
rect 28000 57254 28028 57394
rect 22652 57248 22704 57254
rect 27988 57248 28040 57254
rect 22652 57190 22704 57196
rect 27986 57216 27988 57225
rect 28040 57216 28042 57225
rect 15936 56704 15988 56710
rect 15936 56646 15988 56652
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 2412 22704 2464 22710
rect 2412 22646 2464 22652
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2424 5914 2452 22646
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2424 5710 2452 5850
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 1766 5264 1822 5273
rect 1766 5199 1822 5208
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 12452 2650 12480 26794
rect 15948 22982 15976 56646
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 15936 22976 15988 22982
rect 15936 22918 15988 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 22112 18426 22140 19110
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 22112 17338 22140 18362
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22112 16658 22140 17274
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 22112 16250 22140 16594
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21376 14822 21404 14962
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12452 2446 12480 2586
rect 21376 2514 21404 14758
rect 22204 2582 22232 21422
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22296 18970 22324 19246
rect 22284 18964 22336 18970
rect 22284 18906 22336 18912
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22296 18222 22324 18566
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22572 15570 22600 17138
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22388 14414 22416 15302
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22664 5681 22692 57190
rect 27986 57151 28042 57160
rect 27068 24200 27120 24206
rect 27068 24142 27120 24148
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 22848 22574 22876 23054
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22848 20534 22876 22510
rect 23400 22506 23428 23054
rect 23388 22500 23440 22506
rect 23388 22442 23440 22448
rect 23112 22432 23164 22438
rect 23112 22374 23164 22380
rect 23124 22030 23152 22374
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 24032 22024 24084 22030
rect 24032 21966 24084 21972
rect 23400 21486 23428 21966
rect 23756 21956 23808 21962
rect 23756 21898 23808 21904
rect 23768 21554 23796 21898
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23676 21146 23704 21490
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23860 20942 23888 21830
rect 24044 21622 24072 21966
rect 24032 21616 24084 21622
rect 24032 21558 24084 21564
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 23296 20528 23348 20534
rect 23296 20470 23348 20476
rect 23308 18222 23336 20470
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 23584 20058 23612 20402
rect 23940 20324 23992 20330
rect 23940 20266 23992 20272
rect 23952 20058 23980 20266
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23768 18766 23796 19450
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23860 18630 23888 19246
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23860 18358 23888 18566
rect 23952 18426 23980 19994
rect 24044 19854 24072 20402
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23940 18420 23992 18426
rect 23940 18362 23992 18368
rect 23848 18352 23900 18358
rect 23848 18294 23900 18300
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23308 17882 23336 18158
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23768 17134 23796 17614
rect 23756 17128 23808 17134
rect 23756 17070 23808 17076
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23584 16250 23612 16934
rect 23768 16794 23796 17070
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23768 16250 23796 16594
rect 23860 16522 23888 18294
rect 24044 17882 24072 19790
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 24044 17202 24072 17682
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23584 15706 23612 16186
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23768 15502 23796 16186
rect 23860 16182 23888 16458
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 24032 15632 24084 15638
rect 24032 15574 24084 15580
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 22848 15094 22876 15438
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 22836 15088 22888 15094
rect 22836 15030 22888 15036
rect 23308 14414 23336 15302
rect 23584 15162 23612 15438
rect 24044 15162 24072 15574
rect 24308 15564 24360 15570
rect 24308 15506 24360 15512
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 24320 14958 24348 15506
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 24136 14618 24164 14894
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 23296 14408 23348 14414
rect 23296 14350 23348 14356
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24032 11824 24084 11830
rect 24032 11766 24084 11772
rect 23848 11076 23900 11082
rect 23848 11018 23900 11024
rect 23860 10062 23888 11018
rect 23848 10056 23900 10062
rect 23848 9998 23900 10004
rect 23860 7478 23888 9998
rect 24044 8838 24072 11766
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 24044 8430 24072 8774
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 24136 6458 24164 9590
rect 24320 6934 24348 12786
rect 24412 11626 24440 23598
rect 25056 22506 25084 23666
rect 27080 23118 27108 24142
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 27540 23322 27568 23666
rect 27528 23316 27580 23322
rect 27528 23258 27580 23264
rect 27632 23202 27660 24142
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27816 23730 27844 24006
rect 28736 23866 28764 57462
rect 32232 57458 32260 59200
rect 38028 57594 38056 59200
rect 43180 57594 43208 59200
rect 48976 57594 49004 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 54772 57594 54800 59200
rect 58268 57594 58296 59871
rect 38016 57588 38068 57594
rect 38016 57530 38068 57536
rect 43168 57588 43220 57594
rect 43168 57530 43220 57536
rect 48964 57588 49016 57594
rect 48964 57530 49016 57536
rect 54760 57588 54812 57594
rect 54760 57530 54812 57536
rect 58256 57588 58308 57594
rect 58256 57530 58308 57536
rect 32220 57452 32272 57458
rect 32220 57394 32272 57400
rect 43720 57452 43772 57458
rect 43720 57394 43772 57400
rect 49240 57452 49292 57458
rect 49240 57394 49292 57400
rect 55496 57452 55548 57458
rect 55496 57394 55548 57400
rect 57704 57452 57756 57458
rect 57704 57394 57756 57400
rect 32036 57384 32088 57390
rect 32036 57326 32088 57332
rect 31668 24744 31720 24750
rect 31668 24686 31720 24692
rect 31680 24290 31708 24686
rect 31496 24262 31708 24290
rect 31496 24206 31524 24262
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 31588 23866 31616 24142
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 31576 23860 31628 23866
rect 31576 23802 31628 23808
rect 30564 23792 30616 23798
rect 30564 23734 30616 23740
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 27540 23174 27660 23202
rect 27540 23118 27568 23174
rect 28000 23118 28028 23666
rect 30208 23322 30236 23666
rect 30196 23316 30248 23322
rect 30196 23258 30248 23264
rect 28632 23248 28684 23254
rect 28632 23190 28684 23196
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 26700 23112 26752 23118
rect 26700 23054 26752 23060
rect 27068 23112 27120 23118
rect 27068 23054 27120 23060
rect 27528 23112 27580 23118
rect 27528 23054 27580 23060
rect 27988 23112 28040 23118
rect 27988 23054 28040 23060
rect 26252 22574 26280 23054
rect 26712 22642 26740 23054
rect 27080 22778 27108 23054
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 27540 22658 27568 23054
rect 26700 22636 26752 22642
rect 26700 22578 26752 22584
rect 27448 22630 27568 22658
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 25044 22500 25096 22506
rect 25044 22442 25096 22448
rect 25056 22098 25084 22442
rect 25872 22432 25924 22438
rect 25872 22374 25924 22380
rect 24768 22092 24820 22098
rect 25044 22092 25096 22098
rect 24820 22052 24900 22080
rect 24768 22034 24820 22040
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24492 21888 24544 21894
rect 24492 21830 24544 21836
rect 24504 21690 24532 21830
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24688 21146 24716 21966
rect 24872 21894 24900 22052
rect 25044 22034 25096 22040
rect 25884 22030 25912 22374
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 26424 22024 26476 22030
rect 26424 21966 26476 21972
rect 24860 21888 24912 21894
rect 24860 21830 24912 21836
rect 24872 21690 24900 21830
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24676 21140 24728 21146
rect 24676 21082 24728 21088
rect 24780 20874 24808 21490
rect 24872 20874 24900 21626
rect 24952 21548 25004 21554
rect 24952 21490 25004 21496
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24964 21146 24992 21490
rect 24952 21140 25004 21146
rect 24952 21082 25004 21088
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24780 20602 24808 20810
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 24492 20392 24544 20398
rect 24492 20334 24544 20340
rect 24504 19922 24532 20334
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 25056 19786 25084 21490
rect 25700 21350 25728 21966
rect 26056 21888 26108 21894
rect 26056 21830 26108 21836
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26068 21554 26096 21830
rect 26252 21690 26280 21830
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26056 21548 26108 21554
rect 26056 21490 26108 21496
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25516 20874 25544 21286
rect 25504 20868 25556 20874
rect 25504 20810 25556 20816
rect 25516 20466 25544 20810
rect 25700 20602 25728 21286
rect 26068 21010 26096 21490
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25044 19780 25096 19786
rect 25044 19722 25096 19728
rect 25056 19514 25084 19722
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 25136 19236 25188 19242
rect 25136 19178 25188 19184
rect 25148 18766 25176 19178
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24780 17746 24808 18226
rect 24872 17746 24900 18294
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 24768 17740 24820 17746
rect 24768 17682 24820 17688
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24780 17338 24808 17682
rect 24964 17626 24992 17818
rect 25056 17678 25084 18362
rect 25148 18290 25176 18702
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 24872 17598 24992 17626
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 24872 17202 24900 17598
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24768 16516 24820 16522
rect 24768 16458 24820 16464
rect 24780 15162 24808 16458
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24780 15042 24808 15098
rect 24688 15014 24808 15042
rect 24688 14414 24716 15014
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24492 13184 24544 13190
rect 24492 13126 24544 13132
rect 24504 12782 24532 13126
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24504 12442 24532 12718
rect 24492 12436 24544 12442
rect 24492 12378 24544 12384
rect 24400 11620 24452 11626
rect 24400 11562 24452 11568
rect 24504 10810 24532 12378
rect 24780 11898 24808 14894
rect 24872 13410 24900 17138
rect 25056 16046 25084 17614
rect 25148 17610 25176 18226
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25044 16040 25096 16046
rect 25044 15982 25096 15988
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24964 14346 24992 15642
rect 24952 14340 25004 14346
rect 24952 14282 25004 14288
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 24964 13530 24992 13874
rect 24952 13524 25004 13530
rect 25004 13484 25084 13512
rect 24952 13466 25004 13472
rect 24872 13382 24992 13410
rect 24860 13252 24912 13258
rect 24860 13194 24912 13200
rect 24872 12850 24900 13194
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24964 11898 24992 13382
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 10849 24624 11494
rect 24964 11354 24992 11698
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 25056 11150 25084 13484
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 24582 10840 24638 10849
rect 24492 10804 24544 10810
rect 24582 10775 24638 10784
rect 24492 10746 24544 10752
rect 25240 10742 25268 11766
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24688 10266 24716 10542
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24780 9994 24808 10610
rect 25240 10470 25268 10678
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 24872 10062 24900 10406
rect 25240 10130 25268 10406
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24584 9988 24636 9994
rect 24584 9930 24636 9936
rect 24768 9988 24820 9994
rect 24768 9930 24820 9936
rect 24596 9518 24624 9930
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24964 7410 24992 9318
rect 25240 7886 25268 10066
rect 25332 8634 25360 19790
rect 25516 19514 25544 19858
rect 26068 19514 26096 20946
rect 26148 20936 26200 20942
rect 26252 20890 26280 21626
rect 26436 21554 26464 21966
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26436 20942 26464 21490
rect 26200 20884 26280 20890
rect 26148 20878 26280 20884
rect 26424 20936 26476 20942
rect 26424 20878 26476 20884
rect 26160 20862 26280 20878
rect 26252 20602 26280 20862
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25424 19174 25452 19314
rect 26252 19310 26280 19790
rect 26344 19718 26372 20538
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 26436 19854 26464 20402
rect 26516 20324 26568 20330
rect 26516 20266 26568 20272
rect 26528 19990 26556 20266
rect 26516 19984 26568 19990
rect 26516 19926 26568 19932
rect 26424 19848 26476 19854
rect 26424 19790 26476 19796
rect 26620 19786 26648 20402
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26344 19310 26372 19654
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26332 19304 26384 19310
rect 26332 19246 26384 19252
rect 26516 19304 26568 19310
rect 26620 19292 26648 19722
rect 26568 19264 26648 19292
rect 26516 19246 26568 19252
rect 25412 19168 25464 19174
rect 25412 19110 25464 19116
rect 25424 15706 25452 19110
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 18290 25636 18566
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25516 17338 25544 18226
rect 25700 17610 25728 18634
rect 25792 17882 25820 18702
rect 26252 18426 26280 19246
rect 26344 18426 26372 19246
rect 26424 18692 26476 18698
rect 26424 18634 26476 18640
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 26436 18358 26464 18634
rect 26424 18352 26476 18358
rect 26424 18294 26476 18300
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 26252 17610 26280 18226
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 25608 17218 25636 17478
rect 25516 17190 25636 17218
rect 25516 16522 25544 17190
rect 25700 16998 25728 17546
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25516 16250 25544 16458
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25410 9072 25466 9081
rect 25410 9007 25466 9016
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25332 8090 25360 8434
rect 25320 8084 25372 8090
rect 25320 8026 25372 8032
rect 25424 7970 25452 9007
rect 25332 7942 25452 7970
rect 25228 7880 25280 7886
rect 25228 7822 25280 7828
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24308 6928 24360 6934
rect 24308 6870 24360 6876
rect 24964 6730 24992 7346
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 25148 6798 25176 7142
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 25056 6118 25084 6734
rect 25240 6458 25268 7822
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25332 6322 25360 7942
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25424 7478 25452 7822
rect 25412 7472 25464 7478
rect 25412 7414 25464 7420
rect 25424 6390 25452 7414
rect 25516 6662 25544 14962
rect 25700 13530 25728 16934
rect 26252 16658 26280 16934
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26160 16250 26188 16526
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 26068 15706 26096 16050
rect 26148 16040 26200 16046
rect 26252 15994 26280 16390
rect 26436 16114 26464 17138
rect 26528 16726 26556 19246
rect 26712 18902 26740 22578
rect 26976 22568 27028 22574
rect 26976 22510 27028 22516
rect 26700 18896 26752 18902
rect 26700 18838 26752 18844
rect 26700 17672 26752 17678
rect 26700 17614 26752 17620
rect 26516 16720 26568 16726
rect 26516 16662 26568 16668
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26516 16448 26568 16454
rect 26516 16390 26568 16396
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26200 15988 26280 15994
rect 26148 15982 26280 15988
rect 26332 16040 26384 16046
rect 26332 15982 26384 15988
rect 26160 15966 26280 15982
rect 26344 15910 26372 15982
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 26252 14618 26280 15438
rect 26240 14612 26292 14618
rect 26240 14554 26292 14560
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 13938 26188 14214
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 25792 12442 25820 13874
rect 26240 13864 26292 13870
rect 25976 13802 26188 13818
rect 26240 13806 26292 13812
rect 25964 13796 26188 13802
rect 26016 13790 26188 13796
rect 25964 13738 26016 13744
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 26068 13394 26096 13670
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 25884 12986 25912 13262
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 25976 12850 26004 13262
rect 26068 12850 26096 13330
rect 26160 12986 26188 13790
rect 26252 13530 26280 13806
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26148 12980 26200 12986
rect 26148 12922 26200 12928
rect 25964 12844 26016 12850
rect 25964 12786 26016 12792
rect 26056 12844 26108 12850
rect 26056 12786 26108 12792
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25688 12368 25740 12374
rect 25688 12310 25740 12316
rect 25700 11762 25728 12310
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25700 11286 25728 11698
rect 25688 11280 25740 11286
rect 25688 11222 25740 11228
rect 25688 11008 25740 11014
rect 25688 10950 25740 10956
rect 25700 9926 25728 10950
rect 25688 9920 25740 9926
rect 25688 9862 25740 9868
rect 25700 9042 25728 9862
rect 25792 9654 25820 12378
rect 26056 11756 26108 11762
rect 26056 11698 26108 11704
rect 25872 11688 25924 11694
rect 25872 11630 25924 11636
rect 25780 9648 25832 9654
rect 25780 9590 25832 9596
rect 25688 9036 25740 9042
rect 25688 8978 25740 8984
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25608 8566 25636 8774
rect 25884 8566 25912 11630
rect 26068 11354 26096 11698
rect 26240 11620 26292 11626
rect 26240 11562 26292 11568
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 25964 11144 26016 11150
rect 25964 11086 26016 11092
rect 25976 10062 26004 11086
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 25964 10056 26016 10062
rect 25964 9998 26016 10004
rect 25976 9586 26004 9998
rect 25964 9580 26016 9586
rect 25964 9522 26016 9528
rect 25964 9104 26016 9110
rect 25964 9046 26016 9052
rect 25596 8560 25648 8566
rect 25596 8502 25648 8508
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 25780 8016 25832 8022
rect 25780 7958 25832 7964
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 25412 6384 25464 6390
rect 25412 6326 25464 6332
rect 25320 6316 25372 6322
rect 25320 6258 25372 6264
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 22650 5672 22706 5681
rect 22650 5607 22706 5616
rect 25332 4554 25360 6258
rect 25792 6254 25820 7958
rect 25884 7546 25912 8502
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 25976 7410 26004 9046
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25872 6792 25924 6798
rect 25872 6734 25924 6740
rect 25780 6248 25832 6254
rect 25780 6190 25832 6196
rect 25792 5846 25820 6190
rect 25884 5914 25912 6734
rect 25872 5908 25924 5914
rect 25872 5850 25924 5856
rect 25780 5840 25832 5846
rect 25780 5782 25832 5788
rect 25976 5302 26004 7346
rect 26068 6610 26096 8910
rect 26160 6730 26188 11018
rect 26252 7410 26280 11562
rect 26344 10266 26372 15846
rect 26436 15162 26464 16050
rect 26528 15638 26556 16390
rect 26620 16250 26648 16526
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26516 15632 26568 15638
rect 26516 15574 26568 15580
rect 26424 15156 26476 15162
rect 26424 15098 26476 15104
rect 26528 15094 26556 15574
rect 26516 15088 26568 15094
rect 26516 15030 26568 15036
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26436 12850 26464 13942
rect 26528 13938 26556 14282
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26436 11694 26464 12786
rect 26608 12096 26660 12102
rect 26606 12064 26608 12073
rect 26660 12064 26662 12073
rect 26606 11999 26662 12008
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26516 11620 26568 11626
rect 26516 11562 26568 11568
rect 26424 10736 26476 10742
rect 26424 10678 26476 10684
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26332 9988 26384 9994
rect 26332 9930 26384 9936
rect 26344 9897 26372 9930
rect 26330 9888 26386 9897
rect 26330 9823 26386 9832
rect 26436 9382 26464 10678
rect 26528 10470 26556 11562
rect 26516 10464 26568 10470
rect 26516 10406 26568 10412
rect 26606 10432 26662 10441
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 26528 8906 26556 10406
rect 26606 10367 26662 10376
rect 26620 10062 26648 10367
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26516 8900 26568 8906
rect 26516 8842 26568 8848
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 26344 8430 26372 8774
rect 26620 8566 26648 9454
rect 26712 8634 26740 17614
rect 26988 15978 27016 22510
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 27160 22024 27212 22030
rect 27160 21966 27212 21972
rect 27080 20058 27108 21966
rect 27172 21690 27200 21966
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27448 21622 27476 22630
rect 27528 22568 27580 22574
rect 27528 22510 27580 22516
rect 27540 22234 27568 22510
rect 27528 22228 27580 22234
rect 27528 22170 27580 22176
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27724 21690 27752 21966
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27436 21616 27488 21622
rect 27436 21558 27488 21564
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27724 21010 27752 21422
rect 27896 21140 27948 21146
rect 27896 21082 27948 21088
rect 27712 21004 27764 21010
rect 27712 20946 27764 20952
rect 27528 20324 27580 20330
rect 27528 20266 27580 20272
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 27172 18290 27200 19246
rect 27540 18970 27568 20266
rect 27724 19310 27752 20946
rect 27804 20800 27856 20806
rect 27804 20742 27856 20748
rect 27712 19304 27764 19310
rect 27712 19246 27764 19252
rect 27528 18964 27580 18970
rect 27528 18906 27580 18912
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27252 18216 27304 18222
rect 27252 18158 27304 18164
rect 27264 17814 27292 18158
rect 27540 18086 27568 18906
rect 27528 18080 27580 18086
rect 27528 18022 27580 18028
rect 27816 17882 27844 20742
rect 27908 20466 27936 21082
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27908 18426 27936 20402
rect 28000 19990 28028 23054
rect 28540 23044 28592 23050
rect 28540 22986 28592 22992
rect 28552 22574 28580 22986
rect 28644 22658 28672 23190
rect 30576 23118 30604 23734
rect 31300 23656 31352 23662
rect 31300 23598 31352 23604
rect 31024 23248 31076 23254
rect 31024 23190 31076 23196
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 30564 23112 30616 23118
rect 30564 23054 30616 23060
rect 30748 23112 30800 23118
rect 30748 23054 30800 23060
rect 29012 22778 29040 23054
rect 29460 23044 29512 23050
rect 29460 22986 29512 22992
rect 29000 22772 29052 22778
rect 29000 22714 29052 22720
rect 28644 22642 28856 22658
rect 29472 22642 29500 22986
rect 30288 22976 30340 22982
rect 30288 22918 30340 22924
rect 30300 22642 30328 22918
rect 30576 22642 30604 23054
rect 28644 22636 28868 22642
rect 28644 22630 28816 22636
rect 28540 22568 28592 22574
rect 28540 22510 28592 22516
rect 28644 22234 28672 22630
rect 28816 22578 28868 22584
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30564 22636 30616 22642
rect 30564 22578 30616 22584
rect 28632 22228 28684 22234
rect 28632 22170 28684 22176
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 30012 21548 30064 21554
rect 30012 21490 30064 21496
rect 28092 21146 28120 21490
rect 28632 21344 28684 21350
rect 28632 21286 28684 21292
rect 28080 21140 28132 21146
rect 28080 21082 28132 21088
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28460 20602 28488 20878
rect 28540 20868 28592 20874
rect 28540 20810 28592 20816
rect 28552 20602 28580 20810
rect 28448 20596 28500 20602
rect 28448 20538 28500 20544
rect 28540 20596 28592 20602
rect 28540 20538 28592 20544
rect 28644 20534 28672 21286
rect 30024 20942 30052 21490
rect 30300 21146 30328 22578
rect 30576 21622 30604 22578
rect 30760 22234 30788 23054
rect 31036 22642 31064 23190
rect 31312 22642 31340 23598
rect 31680 23202 31708 24262
rect 31588 23174 31708 23202
rect 31024 22636 31076 22642
rect 31024 22578 31076 22584
rect 31300 22636 31352 22642
rect 31300 22578 31352 22584
rect 30748 22228 30800 22234
rect 30748 22170 30800 22176
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 31300 22024 31352 22030
rect 31300 21966 31352 21972
rect 30564 21616 30616 21622
rect 30564 21558 30616 21564
rect 31128 21554 31156 21966
rect 30472 21548 30524 21554
rect 30472 21490 30524 21496
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 30288 21140 30340 21146
rect 30288 21082 30340 21088
rect 30484 20942 30512 21490
rect 30668 21010 30696 21490
rect 31312 21486 31340 21966
rect 31300 21480 31352 21486
rect 31300 21422 31352 21428
rect 30656 21004 30708 21010
rect 30656 20946 30708 20952
rect 30932 21004 30984 21010
rect 30932 20946 30984 20952
rect 30012 20936 30064 20942
rect 30012 20878 30064 20884
rect 30472 20936 30524 20942
rect 30472 20878 30524 20884
rect 30484 20602 30512 20878
rect 30564 20868 30616 20874
rect 30564 20810 30616 20816
rect 30472 20596 30524 20602
rect 30472 20538 30524 20544
rect 28632 20528 28684 20534
rect 28632 20470 28684 20476
rect 30576 20466 30604 20810
rect 30944 20466 30972 20946
rect 31312 20942 31340 21422
rect 31484 21140 31536 21146
rect 31484 21082 31536 21088
rect 31300 20936 31352 20942
rect 31300 20878 31352 20884
rect 31312 20534 31340 20878
rect 31496 20602 31524 21082
rect 31588 20942 31616 23174
rect 31668 23112 31720 23118
rect 31668 23054 31720 23060
rect 31680 22012 31708 23054
rect 31852 22976 31904 22982
rect 31852 22918 31904 22924
rect 31864 22642 31892 22918
rect 31852 22636 31904 22642
rect 31852 22578 31904 22584
rect 31864 22098 31892 22578
rect 31852 22092 31904 22098
rect 31852 22034 31904 22040
rect 31760 22024 31812 22030
rect 31680 21984 31760 22012
rect 31680 21690 31708 21984
rect 31760 21966 31812 21972
rect 31944 21956 31996 21962
rect 31944 21898 31996 21904
rect 31760 21888 31812 21894
rect 31760 21830 31812 21836
rect 31668 21684 31720 21690
rect 31668 21626 31720 21632
rect 31772 21554 31800 21830
rect 31956 21622 31984 21898
rect 31944 21616 31996 21622
rect 31944 21558 31996 21564
rect 31760 21548 31812 21554
rect 31760 21490 31812 21496
rect 31576 20936 31628 20942
rect 31576 20878 31628 20884
rect 31484 20596 31536 20602
rect 31484 20538 31536 20544
rect 31300 20528 31352 20534
rect 31300 20470 31352 20476
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 30564 20460 30616 20466
rect 30564 20402 30616 20408
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 31392 20460 31444 20466
rect 31392 20402 31444 20408
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 27988 19984 28040 19990
rect 27988 19926 28040 19932
rect 28276 19922 28304 19994
rect 28632 19984 28684 19990
rect 28632 19926 28684 19932
rect 28264 19916 28316 19922
rect 28264 19858 28316 19864
rect 28356 19848 28408 19854
rect 28356 19790 28408 19796
rect 28080 19712 28132 19718
rect 28080 19654 28132 19660
rect 28092 19378 28120 19654
rect 28368 19378 28396 19790
rect 28540 19712 28592 19718
rect 28540 19654 28592 19660
rect 28080 19372 28132 19378
rect 28080 19314 28132 19320
rect 28356 19372 28408 19378
rect 28356 19314 28408 19320
rect 28552 19174 28580 19654
rect 28644 19446 28672 19926
rect 29288 19922 29316 20334
rect 29748 20058 29776 20402
rect 29736 20052 29788 20058
rect 29736 19994 29788 20000
rect 29276 19916 29328 19922
rect 29276 19858 29328 19864
rect 28632 19440 28684 19446
rect 28632 19382 28684 19388
rect 28644 19224 28672 19382
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28920 19224 28948 19314
rect 28644 19196 28948 19224
rect 28540 19168 28592 19174
rect 28540 19110 28592 19116
rect 27896 18420 27948 18426
rect 27896 18362 27948 18368
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 27896 18216 27948 18222
rect 28080 18216 28132 18222
rect 27948 18176 28028 18204
rect 27896 18158 27948 18164
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27804 17876 27856 17882
rect 27804 17818 27856 17824
rect 27252 17808 27304 17814
rect 27252 17750 27304 17756
rect 27540 17746 27568 17818
rect 27528 17740 27580 17746
rect 27528 17682 27580 17688
rect 27540 17649 27568 17682
rect 28000 17678 28028 18176
rect 28080 18158 28132 18164
rect 27988 17672 28040 17678
rect 27526 17640 27582 17649
rect 27988 17614 28040 17620
rect 27526 17575 27582 17584
rect 27712 17332 27764 17338
rect 27712 17274 27764 17280
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27632 16658 27660 16934
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27172 16046 27200 16390
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 26976 15972 27028 15978
rect 26976 15914 27028 15920
rect 26988 15094 27016 15914
rect 27448 15706 27476 16050
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 27068 15428 27120 15434
rect 27068 15370 27120 15376
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 26976 15088 27028 15094
rect 26976 15030 27028 15036
rect 27080 15026 27108 15370
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 26884 13796 26936 13802
rect 26884 13738 26936 13744
rect 26896 13462 26924 13738
rect 26884 13456 26936 13462
rect 26884 13398 26936 13404
rect 26896 13326 26924 13398
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26804 12170 26832 12582
rect 26792 12164 26844 12170
rect 26792 12106 26844 12112
rect 26804 10554 26832 12106
rect 26896 12102 26924 13262
rect 26988 13258 27016 13874
rect 26976 13252 27028 13258
rect 26976 13194 27028 13200
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26884 11008 26936 11014
rect 26882 10976 26884 10985
rect 26936 10976 26938 10985
rect 26882 10911 26938 10920
rect 26988 10606 27016 13194
rect 26976 10600 27028 10606
rect 26804 10526 26924 10554
rect 26976 10542 27028 10548
rect 26792 10464 26844 10470
rect 26792 10406 26844 10412
rect 26804 10266 26832 10406
rect 26792 10260 26844 10266
rect 26792 10202 26844 10208
rect 26896 10146 26924 10526
rect 26896 10118 27016 10146
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 26896 9722 26924 9998
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 26792 9648 26844 9654
rect 26792 9590 26844 9596
rect 26804 8838 26832 9590
rect 26988 8974 27016 10118
rect 26976 8968 27028 8974
rect 26976 8910 27028 8916
rect 26792 8832 26844 8838
rect 26792 8774 26844 8780
rect 26700 8628 26752 8634
rect 26700 8570 26752 8576
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 26240 7404 26292 7410
rect 26240 7346 26292 7352
rect 26332 7404 26384 7410
rect 26332 7346 26384 7352
rect 26252 7206 26280 7346
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 26344 6798 26372 7346
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26148 6724 26200 6730
rect 26148 6666 26200 6672
rect 26068 6582 26188 6610
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 26068 5710 26096 6258
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 26068 5545 26096 5646
rect 26054 5536 26110 5545
rect 26054 5471 26110 5480
rect 25964 5296 26016 5302
rect 25964 5238 26016 5244
rect 26068 4826 26096 5471
rect 26160 5370 26188 6582
rect 26332 6248 26384 6254
rect 26332 6190 26384 6196
rect 26148 5364 26200 5370
rect 26148 5306 26200 5312
rect 26344 5234 26372 6190
rect 26436 5642 26464 8298
rect 26804 7954 26832 8774
rect 26884 8288 26936 8294
rect 26884 8230 26936 8236
rect 26896 7954 26924 8230
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26884 7948 26936 7954
rect 26884 7890 26936 7896
rect 26528 6610 26556 7890
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 26988 7478 27016 7822
rect 27080 7546 27108 14962
rect 27540 14822 27568 15370
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27632 14618 27660 14962
rect 27620 14612 27672 14618
rect 27620 14554 27672 14560
rect 27724 14482 27752 17274
rect 28000 16726 28028 17614
rect 28092 17542 28120 18158
rect 28184 17678 28212 18226
rect 28552 18086 28580 19110
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28540 18080 28592 18086
rect 28540 18022 28592 18028
rect 28276 17678 28304 18022
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 28264 17672 28316 17678
rect 28264 17614 28316 17620
rect 28080 17536 28132 17542
rect 28080 17478 28132 17484
rect 28184 17490 28212 17614
rect 28264 17536 28316 17542
rect 28184 17484 28264 17490
rect 28184 17478 28316 17484
rect 28184 17462 28304 17478
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 27988 16720 28040 16726
rect 27988 16662 28040 16668
rect 27896 15972 27948 15978
rect 27896 15914 27948 15920
rect 27908 15638 27936 15914
rect 28092 15706 28120 17138
rect 28448 16992 28500 16998
rect 28448 16934 28500 16940
rect 28460 16522 28488 16934
rect 28448 16516 28500 16522
rect 28448 16458 28500 16464
rect 28460 15910 28488 16458
rect 28448 15904 28500 15910
rect 28448 15846 28500 15852
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 27896 15632 27948 15638
rect 27896 15574 27948 15580
rect 27908 14498 27936 15574
rect 27988 15496 28040 15502
rect 27988 15438 28040 15444
rect 28000 15026 28028 15438
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27816 14470 27936 14498
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27172 11830 27200 12786
rect 27252 12708 27304 12714
rect 27252 12650 27304 12656
rect 27344 12708 27396 12714
rect 27344 12650 27396 12656
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 27160 11688 27212 11694
rect 27160 11630 27212 11636
rect 27172 10130 27200 11630
rect 27264 11558 27292 12650
rect 27356 12306 27384 12650
rect 27448 12442 27476 12786
rect 27632 12730 27660 14350
rect 27816 13462 27844 14470
rect 27896 14272 27948 14278
rect 27896 14214 27948 14220
rect 27908 14006 27936 14214
rect 27896 14000 27948 14006
rect 27896 13942 27948 13948
rect 27804 13456 27856 13462
rect 27804 13398 27856 13404
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27724 12850 27752 13126
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27632 12702 27752 12730
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27448 12306 27660 12322
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 27436 12300 27660 12306
rect 27488 12294 27660 12300
rect 27436 12242 27488 12248
rect 27528 12232 27580 12238
rect 27528 12174 27580 12180
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27448 11354 27476 11698
rect 27540 11694 27568 12174
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27528 11552 27580 11558
rect 27632 11506 27660 12294
rect 27580 11500 27660 11506
rect 27528 11494 27660 11500
rect 27540 11478 27660 11494
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27344 11280 27396 11286
rect 27344 11222 27396 11228
rect 27252 11008 27304 11014
rect 27252 10950 27304 10956
rect 27264 10470 27292 10950
rect 27356 10674 27384 11222
rect 27436 10736 27488 10742
rect 27436 10678 27488 10684
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27344 10532 27396 10538
rect 27344 10474 27396 10480
rect 27252 10464 27304 10470
rect 27252 10406 27304 10412
rect 27160 10124 27212 10130
rect 27160 10066 27212 10072
rect 27264 9654 27292 10406
rect 27356 10062 27384 10474
rect 27448 10169 27476 10678
rect 27434 10160 27490 10169
rect 27434 10095 27490 10104
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 27540 9874 27568 11478
rect 27618 11112 27674 11121
rect 27618 11047 27620 11056
rect 27672 11047 27674 11056
rect 27620 11018 27672 11024
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27356 9846 27568 9874
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 27252 9376 27304 9382
rect 27252 9318 27304 9324
rect 27264 8906 27292 9318
rect 27252 8900 27304 8906
rect 27252 8842 27304 8848
rect 27160 8492 27212 8498
rect 27160 8434 27212 8440
rect 27068 7540 27120 7546
rect 27068 7482 27120 7488
rect 26976 7472 27028 7478
rect 26976 7414 27028 7420
rect 26700 7336 26752 7342
rect 26700 7278 26752 7284
rect 26976 7336 27028 7342
rect 26976 7278 27028 7284
rect 26712 6984 26740 7278
rect 26712 6956 26924 6984
rect 26712 6798 26740 6956
rect 26790 6896 26846 6905
rect 26790 6831 26846 6840
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26804 6730 26832 6831
rect 26792 6724 26844 6730
rect 26792 6666 26844 6672
rect 26528 6582 26740 6610
rect 26712 6254 26740 6582
rect 26700 6248 26752 6254
rect 26700 6190 26752 6196
rect 26424 5636 26476 5642
rect 26424 5578 26476 5584
rect 26332 5228 26384 5234
rect 26332 5170 26384 5176
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26344 4758 26372 5170
rect 26332 4752 26384 4758
rect 26332 4694 26384 4700
rect 25320 4548 25372 4554
rect 25320 4490 25372 4496
rect 26436 3194 26464 5578
rect 26804 5234 26832 6666
rect 26792 5228 26844 5234
rect 26792 5170 26844 5176
rect 26896 5030 26924 6956
rect 26988 5166 27016 7278
rect 27066 7032 27122 7041
rect 27066 6967 27122 6976
rect 27080 6934 27108 6967
rect 27068 6928 27120 6934
rect 27068 6870 27120 6876
rect 27172 5914 27200 8434
rect 27252 8016 27304 8022
rect 27252 7958 27304 7964
rect 27264 6934 27292 7958
rect 27252 6928 27304 6934
rect 27252 6870 27304 6876
rect 27252 6724 27304 6730
rect 27356 6712 27384 9846
rect 27632 9761 27660 10610
rect 27724 10266 27752 12702
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27618 9752 27674 9761
rect 27618 9687 27674 9696
rect 27632 9518 27660 9687
rect 27816 9654 27844 13262
rect 27896 12980 27948 12986
rect 27896 12922 27948 12928
rect 27908 11898 27936 12922
rect 28000 12782 28028 14962
rect 28092 12918 28120 15642
rect 28264 14816 28316 14822
rect 28264 14758 28316 14764
rect 28276 14482 28304 14758
rect 28172 14476 28224 14482
rect 28172 14418 28224 14424
rect 28264 14476 28316 14482
rect 28264 14418 28316 14424
rect 28080 12912 28132 12918
rect 28080 12854 28132 12860
rect 28184 12850 28212 14418
rect 28276 14346 28304 14418
rect 28264 14340 28316 14346
rect 28264 14282 28316 14288
rect 28172 12844 28224 12850
rect 28172 12786 28224 12792
rect 27988 12776 28040 12782
rect 27988 12718 28040 12724
rect 28080 12164 28132 12170
rect 28080 12106 28132 12112
rect 27896 11892 27948 11898
rect 27896 11834 27948 11840
rect 28092 11830 28120 12106
rect 28080 11824 28132 11830
rect 28080 11766 28132 11772
rect 27896 11212 27948 11218
rect 27896 11154 27948 11160
rect 27804 9648 27856 9654
rect 27804 9590 27856 9596
rect 27620 9512 27672 9518
rect 27620 9454 27672 9460
rect 27712 9376 27764 9382
rect 27712 9318 27764 9324
rect 27620 8968 27672 8974
rect 27618 8936 27620 8945
rect 27672 8936 27674 8945
rect 27724 8922 27752 9318
rect 27816 9110 27844 9590
rect 27908 9586 27936 11154
rect 28184 11150 28212 12786
rect 28354 12200 28410 12209
rect 28354 12135 28356 12144
rect 28408 12135 28410 12144
rect 28356 12106 28408 12112
rect 28264 11756 28316 11762
rect 28264 11698 28316 11704
rect 28276 11354 28304 11698
rect 28264 11348 28316 11354
rect 28264 11290 28316 11296
rect 28368 11150 28396 12106
rect 28172 11144 28224 11150
rect 28172 11086 28224 11092
rect 28356 11144 28408 11150
rect 28356 11086 28408 11092
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 28276 10985 28304 11018
rect 28262 10976 28318 10985
rect 28262 10911 28318 10920
rect 28080 10464 28132 10470
rect 28460 10418 28488 15846
rect 28540 15496 28592 15502
rect 28540 15438 28592 15444
rect 28552 14618 28580 15438
rect 28644 15366 28672 19196
rect 29288 18766 29316 19858
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29552 19780 29604 19786
rect 29552 19722 29604 19728
rect 29564 19242 29592 19722
rect 29932 19378 29960 19790
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 30380 19372 30432 19378
rect 30380 19314 30432 19320
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29552 19236 29604 19242
rect 29552 19178 29604 19184
rect 29276 18760 29328 18766
rect 29276 18702 29328 18708
rect 29092 18692 29144 18698
rect 29092 18634 29144 18640
rect 28908 18080 28960 18086
rect 28960 18028 29040 18034
rect 28908 18022 29040 18028
rect 28920 18006 29040 18022
rect 29012 17066 29040 18006
rect 29104 17746 29132 18634
rect 29092 17740 29144 17746
rect 29092 17682 29144 17688
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 29000 17060 29052 17066
rect 29000 17002 29052 17008
rect 29012 16794 29040 17002
rect 29000 16788 29052 16794
rect 29000 16730 29052 16736
rect 29012 16250 29040 16730
rect 29104 16522 29132 17138
rect 29092 16516 29144 16522
rect 29092 16458 29144 16464
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 28816 15632 28868 15638
rect 28816 15574 28868 15580
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28632 15360 28684 15366
rect 28736 15337 28764 15438
rect 28632 15302 28684 15308
rect 28722 15328 28778 15337
rect 28722 15263 28778 15272
rect 28828 15026 28856 15574
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 28908 15360 28960 15366
rect 28908 15302 28960 15308
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 28540 14612 28592 14618
rect 28540 14554 28592 14560
rect 28552 11762 28580 14554
rect 28722 14104 28778 14113
rect 28722 14039 28724 14048
rect 28776 14039 28778 14048
rect 28724 14010 28776 14016
rect 28736 13870 28764 14010
rect 28828 13938 28856 14962
rect 28920 14890 28948 15302
rect 29012 15162 29040 15438
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 28908 14884 28960 14890
rect 28908 14826 28960 14832
rect 29104 14550 29132 16458
rect 29184 14952 29236 14958
rect 29184 14894 29236 14900
rect 29092 14544 29144 14550
rect 29092 14486 29144 14492
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28724 12640 28776 12646
rect 28724 12582 28776 12588
rect 28736 12238 28764 12582
rect 28828 12374 28856 13874
rect 28920 13802 28948 14214
rect 28908 13796 28960 13802
rect 28908 13738 28960 13744
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28920 12986 28948 13262
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 28816 12368 28868 12374
rect 28816 12310 28868 12316
rect 28724 12232 28776 12238
rect 28724 12174 28776 12180
rect 28632 12096 28684 12102
rect 28632 12038 28684 12044
rect 28540 11756 28592 11762
rect 28540 11698 28592 11704
rect 28552 10470 28580 11698
rect 28644 10742 28672 12038
rect 28724 11688 28776 11694
rect 28724 11630 28776 11636
rect 28632 10736 28684 10742
rect 28632 10678 28684 10684
rect 28540 10464 28592 10470
rect 28080 10406 28132 10412
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 27896 9580 27948 9586
rect 27896 9522 27948 9528
rect 27804 9104 27856 9110
rect 27804 9046 27856 9052
rect 27908 8974 27936 9522
rect 27896 8968 27948 8974
rect 27724 8894 27844 8922
rect 27896 8910 27948 8916
rect 27618 8871 27674 8880
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27448 8090 27476 8366
rect 27816 8090 27844 8894
rect 27894 8800 27950 8809
rect 27894 8735 27950 8744
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 27528 7812 27580 7818
rect 27528 7754 27580 7760
rect 27436 7268 27488 7274
rect 27436 7210 27488 7216
rect 27448 7002 27476 7210
rect 27436 6996 27488 7002
rect 27436 6938 27488 6944
rect 27540 6798 27568 7754
rect 27618 7440 27674 7449
rect 27618 7375 27620 7384
rect 27672 7375 27674 7384
rect 27620 7346 27672 7352
rect 27632 7188 27660 7346
rect 27712 7200 27764 7206
rect 27632 7160 27712 7188
rect 27712 7142 27764 7148
rect 27620 6996 27672 7002
rect 27620 6938 27672 6944
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27304 6684 27384 6712
rect 27252 6666 27304 6672
rect 27356 6225 27384 6684
rect 27448 6254 27476 6734
rect 27436 6248 27488 6254
rect 27342 6216 27398 6225
rect 27436 6190 27488 6196
rect 27342 6151 27398 6160
rect 27160 5908 27212 5914
rect 27160 5850 27212 5856
rect 27356 5710 27384 6151
rect 27632 5778 27660 6938
rect 27816 6730 27844 8026
rect 27908 7342 27936 8735
rect 28000 7449 28028 10202
rect 28092 10062 28120 10406
rect 28184 10390 28488 10418
rect 28538 10432 28540 10441
rect 28592 10432 28594 10441
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 28078 9888 28134 9897
rect 28078 9823 28134 9832
rect 27986 7440 28042 7449
rect 27986 7375 28042 7384
rect 27896 7336 27948 7342
rect 27988 7336 28040 7342
rect 27896 7278 27948 7284
rect 27986 7304 27988 7313
rect 28040 7304 28042 7313
rect 27986 7239 28042 7248
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27620 5772 27672 5778
rect 27620 5714 27672 5720
rect 27344 5704 27396 5710
rect 27264 5664 27344 5692
rect 26976 5160 27028 5166
rect 26976 5102 27028 5108
rect 26884 5024 26936 5030
rect 26884 4966 26936 4972
rect 27264 4826 27292 5664
rect 27344 5646 27396 5652
rect 27344 5568 27396 5574
rect 27344 5510 27396 5516
rect 27356 5370 27384 5510
rect 27632 5409 27660 5714
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27618 5400 27674 5409
rect 27344 5364 27396 5370
rect 27618 5335 27674 5344
rect 27344 5306 27396 5312
rect 27724 4826 27752 5646
rect 27816 5234 27844 6666
rect 28000 6338 28028 7239
rect 28092 6866 28120 9823
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 27908 6310 28028 6338
rect 28080 6384 28132 6390
rect 28080 6326 28132 6332
rect 27908 6118 27936 6310
rect 27896 6112 27948 6118
rect 27896 6054 27948 6060
rect 27988 6112 28040 6118
rect 27988 6054 28040 6060
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27252 4820 27304 4826
rect 27252 4762 27304 4768
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27816 4010 27844 4626
rect 27804 4004 27856 4010
rect 27804 3946 27856 3952
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 27908 2990 27936 6054
rect 28000 5098 28028 6054
rect 27988 5092 28040 5098
rect 27988 5034 28040 5040
rect 28092 4622 28120 6326
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 28092 4146 28120 4558
rect 28184 4486 28212 10390
rect 28538 10367 28594 10376
rect 28446 10296 28502 10305
rect 28644 10266 28672 10678
rect 28446 10231 28448 10240
rect 28500 10231 28502 10240
rect 28632 10260 28684 10266
rect 28448 10202 28500 10208
rect 28632 10202 28684 10208
rect 28540 10192 28592 10198
rect 28262 10160 28318 10169
rect 28540 10134 28592 10140
rect 28262 10095 28318 10104
rect 28276 9586 28304 10095
rect 28356 9920 28408 9926
rect 28356 9862 28408 9868
rect 28368 9654 28396 9862
rect 28552 9654 28580 10134
rect 28356 9648 28408 9654
rect 28356 9590 28408 9596
rect 28540 9648 28592 9654
rect 28540 9590 28592 9596
rect 28264 9580 28316 9586
rect 28264 9522 28316 9528
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 28264 9104 28316 9110
rect 28262 9072 28264 9081
rect 28316 9072 28318 9081
rect 28262 9007 28318 9016
rect 28264 8560 28316 8566
rect 28264 8502 28316 8508
rect 28276 7750 28304 8502
rect 28368 8362 28396 9318
rect 28448 8900 28500 8906
rect 28448 8842 28500 8848
rect 28460 8498 28488 8842
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 28356 8356 28408 8362
rect 28552 8344 28580 9590
rect 28632 9580 28684 9586
rect 28632 9522 28684 9528
rect 28644 8634 28672 9522
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28632 8492 28684 8498
rect 28632 8434 28684 8440
rect 28356 8298 28408 8304
rect 28460 8316 28580 8344
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28276 5098 28304 7686
rect 28460 7342 28488 8316
rect 28540 7880 28592 7886
rect 28644 7868 28672 8434
rect 28592 7840 28672 7868
rect 28540 7822 28592 7828
rect 28448 7336 28500 7342
rect 28448 7278 28500 7284
rect 28354 7032 28410 7041
rect 28354 6967 28356 6976
rect 28408 6967 28410 6976
rect 28356 6938 28408 6944
rect 28552 6866 28580 7822
rect 28736 7478 28764 11630
rect 29012 11354 29040 13262
rect 29104 12850 29132 13330
rect 29196 13190 29224 14894
rect 29184 13184 29236 13190
rect 29184 13126 29236 13132
rect 29196 12986 29224 13126
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 29092 12844 29144 12850
rect 29092 12786 29144 12792
rect 28816 11348 28868 11354
rect 28816 11290 28868 11296
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 28828 10606 28856 11290
rect 28908 11280 28960 11286
rect 28960 11228 29040 11234
rect 28908 11222 29040 11228
rect 28920 11206 29040 11222
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28920 10985 28948 11086
rect 28906 10976 28962 10985
rect 28906 10911 28962 10920
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28908 10260 28960 10266
rect 28908 10202 28960 10208
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 28828 9722 28856 9998
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 28816 9512 28868 9518
rect 28816 9454 28868 9460
rect 28828 8022 28856 9454
rect 28920 9217 28948 10202
rect 28906 9208 28962 9217
rect 28906 9143 28962 9152
rect 28920 9110 28948 9143
rect 28908 9104 28960 9110
rect 28908 9046 28960 9052
rect 29012 8974 29040 11206
rect 29104 10062 29132 12786
rect 29288 12434 29316 18702
rect 29564 18290 29592 19178
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29656 18154 29684 19246
rect 29840 18970 29868 19246
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 29840 18154 29868 18906
rect 29932 18290 29960 19314
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 30024 18426 30052 18770
rect 30392 18766 30420 19314
rect 30576 18970 30604 20402
rect 30944 19718 30972 20402
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30564 18964 30616 18970
rect 30564 18906 30616 18912
rect 30380 18760 30432 18766
rect 30380 18702 30432 18708
rect 30012 18420 30064 18426
rect 30012 18362 30064 18368
rect 29920 18284 29972 18290
rect 29920 18226 29972 18232
rect 29644 18148 29696 18154
rect 29644 18090 29696 18096
rect 29828 18148 29880 18154
rect 29828 18090 29880 18096
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29472 16590 29500 16934
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 29472 15910 29500 16526
rect 29460 15904 29512 15910
rect 29460 15846 29512 15852
rect 29656 15162 29684 18090
rect 30288 17264 30340 17270
rect 30288 17206 30340 17212
rect 30300 16726 30328 17206
rect 29736 16720 29788 16726
rect 29736 16662 29788 16668
rect 30288 16720 30340 16726
rect 30288 16662 30340 16668
rect 29748 16114 29776 16662
rect 30196 16584 30248 16590
rect 30196 16526 30248 16532
rect 30208 16114 30236 16526
rect 30300 16454 30328 16662
rect 30288 16448 30340 16454
rect 30288 16390 30340 16396
rect 29736 16108 29788 16114
rect 29736 16050 29788 16056
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 29932 15638 29960 16050
rect 29920 15632 29972 15638
rect 29920 15574 29972 15580
rect 29828 15564 29880 15570
rect 29828 15506 29880 15512
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 29552 14340 29604 14346
rect 29552 14282 29604 14288
rect 29564 13938 29592 14282
rect 29736 14000 29788 14006
rect 29736 13942 29788 13948
rect 29368 13932 29420 13938
rect 29368 13874 29420 13880
rect 29552 13932 29604 13938
rect 29552 13874 29604 13880
rect 29380 13326 29408 13874
rect 29460 13728 29512 13734
rect 29460 13670 29512 13676
rect 29368 13320 29420 13326
rect 29368 13262 29420 13268
rect 29472 12850 29500 13670
rect 29748 13138 29776 13942
rect 29840 13326 29868 15506
rect 29932 15094 29960 15574
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 29920 15088 29972 15094
rect 29920 15030 29972 15036
rect 30012 15020 30064 15026
rect 30012 14962 30064 14968
rect 30104 15020 30156 15026
rect 30104 14962 30156 14968
rect 29920 14612 29972 14618
rect 29920 14554 29972 14560
rect 29932 13938 29960 14554
rect 30024 14074 30052 14962
rect 30012 14068 30064 14074
rect 30012 14010 30064 14016
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 30116 13716 30144 14962
rect 30208 14822 30236 15438
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 30208 13954 30236 14758
rect 30392 14074 30420 18702
rect 31116 18420 31168 18426
rect 31116 18362 31168 18368
rect 31128 18290 31156 18362
rect 30472 18284 30524 18290
rect 30472 18226 30524 18232
rect 31116 18284 31168 18290
rect 31116 18226 31168 18232
rect 30484 17134 30512 18226
rect 31404 17814 31432 20402
rect 31496 20398 31524 20538
rect 31668 20460 31720 20466
rect 31668 20402 31720 20408
rect 31760 20460 31812 20466
rect 31760 20402 31812 20408
rect 31484 20392 31536 20398
rect 31484 20334 31536 20340
rect 31680 20058 31708 20402
rect 31668 20052 31720 20058
rect 31668 19994 31720 20000
rect 31576 19848 31628 19854
rect 31576 19790 31628 19796
rect 31588 19378 31616 19790
rect 31576 19372 31628 19378
rect 31576 19314 31628 19320
rect 31588 18970 31616 19314
rect 31772 19242 31800 20402
rect 31852 19304 31904 19310
rect 31852 19246 31904 19252
rect 31760 19236 31812 19242
rect 31760 19178 31812 19184
rect 31576 18964 31628 18970
rect 31576 18906 31628 18912
rect 31864 18222 31892 19246
rect 31852 18216 31904 18222
rect 31852 18158 31904 18164
rect 31392 17808 31444 17814
rect 31392 17750 31444 17756
rect 31208 17740 31260 17746
rect 31208 17682 31260 17688
rect 30932 17672 30984 17678
rect 30932 17614 30984 17620
rect 30944 17218 30972 17614
rect 31220 17338 31248 17682
rect 31208 17332 31260 17338
rect 31208 17274 31260 17280
rect 30944 17202 31064 17218
rect 30564 17196 30616 17202
rect 30564 17138 30616 17144
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30944 17196 31076 17202
rect 30944 17190 31024 17196
rect 30472 17128 30524 17134
rect 30472 17070 30524 17076
rect 30576 17066 30604 17138
rect 30564 17060 30616 17066
rect 30564 17002 30616 17008
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30484 16182 30512 16526
rect 30576 16250 30604 17002
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30380 14068 30432 14074
rect 30380 14010 30432 14016
rect 30208 13926 30512 13954
rect 30024 13688 30144 13716
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29656 13110 29776 13138
rect 29460 12844 29512 12850
rect 29460 12786 29512 12792
rect 29196 12406 29316 12434
rect 29196 11898 29224 12406
rect 29276 12096 29328 12102
rect 29276 12038 29328 12044
rect 29184 11892 29236 11898
rect 29184 11834 29236 11840
rect 29288 11762 29316 12038
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 29472 11286 29500 12786
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29460 11280 29512 11286
rect 29460 11222 29512 11228
rect 29460 11076 29512 11082
rect 29460 11018 29512 11024
rect 29472 10810 29500 11018
rect 29460 10804 29512 10810
rect 29460 10746 29512 10752
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 29196 10266 29224 10610
rect 29274 10568 29330 10577
rect 29274 10503 29276 10512
rect 29328 10503 29330 10512
rect 29276 10474 29328 10480
rect 29184 10260 29236 10266
rect 29184 10202 29236 10208
rect 29092 10056 29144 10062
rect 29092 9998 29144 10004
rect 29104 9081 29132 9998
rect 29182 9616 29238 9625
rect 29182 9551 29238 9560
rect 29090 9072 29146 9081
rect 29090 9007 29146 9016
rect 29104 8974 29132 9007
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 29092 8968 29144 8974
rect 29092 8910 29144 8916
rect 28816 8016 28868 8022
rect 28816 7958 28868 7964
rect 28908 7812 28960 7818
rect 28908 7754 28960 7760
rect 28724 7472 28776 7478
rect 28724 7414 28776 7420
rect 28920 7342 28948 7754
rect 29012 7750 29040 8910
rect 29196 8362 29224 9551
rect 29368 9444 29420 9450
rect 29368 9386 29420 9392
rect 29380 9110 29408 9386
rect 29368 9104 29420 9110
rect 29368 9046 29420 9052
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29184 8356 29236 8362
rect 29184 8298 29236 8304
rect 29090 7984 29146 7993
rect 29090 7919 29146 7928
rect 29104 7886 29132 7919
rect 29092 7880 29144 7886
rect 29092 7822 29144 7828
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29012 7392 29040 7686
rect 29092 7404 29144 7410
rect 29012 7364 29092 7392
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 28816 6928 28868 6934
rect 28816 6870 28868 6876
rect 28540 6860 28592 6866
rect 28540 6802 28592 6808
rect 28356 6792 28408 6798
rect 28356 6734 28408 6740
rect 28448 6792 28500 6798
rect 28448 6734 28500 6740
rect 28368 6390 28396 6734
rect 28356 6384 28408 6390
rect 28356 6326 28408 6332
rect 28356 6248 28408 6254
rect 28356 6190 28408 6196
rect 28368 5574 28396 6190
rect 28460 6118 28488 6734
rect 28448 6112 28500 6118
rect 28448 6054 28500 6060
rect 28552 5930 28580 6802
rect 28828 6186 28856 6870
rect 29012 6458 29040 7364
rect 29092 7346 29144 7352
rect 29196 6905 29224 8298
rect 29288 8294 29316 8434
rect 29472 8401 29500 10746
rect 29564 9926 29592 12718
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29564 8906 29592 9522
rect 29656 9450 29684 13110
rect 29840 12850 29868 13262
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 29840 12434 29868 12786
rect 29748 12406 29868 12434
rect 29644 9444 29696 9450
rect 29644 9386 29696 9392
rect 29644 8968 29696 8974
rect 29642 8936 29644 8945
rect 29696 8936 29698 8945
rect 29552 8900 29604 8906
rect 29642 8871 29698 8880
rect 29552 8842 29604 8848
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29458 8392 29514 8401
rect 29458 8327 29514 8336
rect 29276 8288 29328 8294
rect 29276 8230 29328 8236
rect 29182 6896 29238 6905
rect 29182 6831 29238 6840
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 28816 6180 28868 6186
rect 28816 6122 28868 6128
rect 28722 6080 28778 6089
rect 28722 6015 28778 6024
rect 28460 5902 28580 5930
rect 28736 5914 28764 6015
rect 28724 5908 28776 5914
rect 28356 5568 28408 5574
rect 28460 5545 28488 5902
rect 28724 5850 28776 5856
rect 28632 5840 28684 5846
rect 28632 5782 28684 5788
rect 28644 5710 28672 5782
rect 28632 5704 28684 5710
rect 28632 5646 28684 5652
rect 29012 5658 29040 6394
rect 29288 6089 29316 8230
rect 29564 7970 29592 8434
rect 29380 7942 29592 7970
rect 29274 6080 29330 6089
rect 29274 6015 29330 6024
rect 28540 5636 28592 5642
rect 28540 5578 28592 5584
rect 28356 5510 28408 5516
rect 28446 5536 28502 5545
rect 28446 5471 28502 5480
rect 28552 5137 28580 5578
rect 28538 5128 28594 5137
rect 28264 5092 28316 5098
rect 28538 5063 28594 5072
rect 28264 5034 28316 5040
rect 28276 4622 28304 5034
rect 28644 5001 28672 5646
rect 29012 5630 29224 5658
rect 28724 5568 28776 5574
rect 28724 5510 28776 5516
rect 28906 5536 28962 5545
rect 28736 5409 28764 5510
rect 28962 5494 29132 5522
rect 28906 5471 28962 5480
rect 28722 5400 28778 5409
rect 28722 5335 28778 5344
rect 28816 5364 28868 5370
rect 28816 5306 28868 5312
rect 28630 4992 28686 5001
rect 28630 4927 28686 4936
rect 28828 4758 28856 5306
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 28816 4752 28868 4758
rect 28816 4694 28868 4700
rect 28356 4684 28408 4690
rect 28356 4626 28408 4632
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28172 4480 28224 4486
rect 28172 4422 28224 4428
rect 28368 4146 28396 4626
rect 28448 4616 28500 4622
rect 28448 4558 28500 4564
rect 28460 4282 28488 4558
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 28080 4140 28132 4146
rect 28080 4082 28132 4088
rect 28356 4140 28408 4146
rect 28356 4082 28408 4088
rect 27988 4072 28040 4078
rect 27986 4040 27988 4049
rect 28040 4040 28042 4049
rect 27986 3975 28042 3984
rect 28460 3738 28488 4218
rect 28448 3732 28500 3738
rect 28448 3674 28500 3680
rect 27896 2984 27948 2990
rect 27896 2926 27948 2932
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 21364 2508 21416 2514
rect 21364 2450 21416 2456
rect 28920 2446 28948 4966
rect 29104 4622 29132 5494
rect 29196 5166 29224 5630
rect 29380 5234 29408 7942
rect 29552 7880 29604 7886
rect 29552 7822 29604 7828
rect 29458 7712 29514 7721
rect 29458 7647 29514 7656
rect 29472 7410 29500 7647
rect 29460 7404 29512 7410
rect 29460 7346 29512 7352
rect 29368 5228 29420 5234
rect 29368 5170 29420 5176
rect 29184 5160 29236 5166
rect 29184 5102 29236 5108
rect 29380 4826 29408 5170
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 29092 4616 29144 4622
rect 29092 4558 29144 4564
rect 29104 4214 29132 4558
rect 29092 4208 29144 4214
rect 29092 4150 29144 4156
rect 29472 4010 29500 7346
rect 29564 5846 29592 7822
rect 29656 7410 29684 8871
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29656 6934 29684 7346
rect 29644 6928 29696 6934
rect 29644 6870 29696 6876
rect 29644 6792 29696 6798
rect 29644 6734 29696 6740
rect 29656 6458 29684 6734
rect 29644 6452 29696 6458
rect 29644 6394 29696 6400
rect 29552 5840 29604 5846
rect 29552 5782 29604 5788
rect 29656 5710 29684 6394
rect 29644 5704 29696 5710
rect 29644 5646 29696 5652
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29564 5234 29592 5510
rect 29552 5228 29604 5234
rect 29552 5170 29604 5176
rect 29460 4004 29512 4010
rect 29460 3946 29512 3952
rect 29748 3738 29776 12406
rect 30024 12170 30052 13688
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 30012 12164 30064 12170
rect 30012 12106 30064 12112
rect 29828 11552 29880 11558
rect 29828 11494 29880 11500
rect 29840 11082 29868 11494
rect 29920 11144 29972 11150
rect 29920 11086 29972 11092
rect 29828 11076 29880 11082
rect 29828 11018 29880 11024
rect 29932 10810 29960 11086
rect 29920 10804 29972 10810
rect 29920 10746 29972 10752
rect 30116 10674 30144 12786
rect 30380 12640 30432 12646
rect 30380 12582 30432 12588
rect 30392 12374 30420 12582
rect 30380 12368 30432 12374
rect 30380 12310 30432 12316
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30288 12232 30340 12238
rect 30288 12174 30340 12180
rect 30208 11257 30236 12174
rect 30300 11801 30328 12174
rect 30380 12164 30432 12170
rect 30380 12106 30432 12112
rect 30286 11792 30342 11801
rect 30286 11727 30342 11736
rect 30194 11248 30250 11257
rect 30300 11218 30328 11727
rect 30392 11393 30420 12106
rect 30378 11384 30434 11393
rect 30378 11319 30434 11328
rect 30194 11183 30250 11192
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 30286 10840 30342 10849
rect 30392 10810 30420 11319
rect 30286 10775 30288 10784
rect 30340 10775 30342 10784
rect 30380 10804 30432 10810
rect 30288 10746 30340 10752
rect 30380 10746 30432 10752
rect 29920 10668 29972 10674
rect 29920 10610 29972 10616
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 29828 10260 29880 10266
rect 29828 10202 29880 10208
rect 29840 10062 29868 10202
rect 29932 10169 29960 10610
rect 30116 10577 30144 10610
rect 30196 10600 30248 10606
rect 30102 10568 30158 10577
rect 30196 10542 30248 10548
rect 30102 10503 30158 10512
rect 30208 10266 30236 10542
rect 30196 10260 30248 10266
rect 30196 10202 30248 10208
rect 29918 10160 29974 10169
rect 29918 10095 29974 10104
rect 29828 10056 29880 10062
rect 29828 9998 29880 10004
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 30116 9926 30144 9998
rect 29920 9920 29972 9926
rect 29920 9862 29972 9868
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 29826 9616 29882 9625
rect 29826 9551 29828 9560
rect 29880 9551 29882 9560
rect 29828 9522 29880 9528
rect 29828 9036 29880 9042
rect 29828 8978 29880 8984
rect 29840 8945 29868 8978
rect 29826 8936 29882 8945
rect 29826 8871 29882 8880
rect 29932 8294 29960 9862
rect 30116 9586 30144 9862
rect 30104 9580 30156 9586
rect 30104 9522 30156 9528
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 30024 9217 30052 9454
rect 30116 9450 30144 9522
rect 30104 9444 30156 9450
rect 30104 9386 30156 9392
rect 30010 9208 30066 9217
rect 30010 9143 30066 9152
rect 30288 9104 30340 9110
rect 30010 9072 30066 9081
rect 30288 9046 30340 9052
rect 30010 9007 30012 9016
rect 30064 9007 30066 9016
rect 30012 8978 30064 8984
rect 30024 8498 30052 8978
rect 30300 8673 30328 9046
rect 30380 8968 30432 8974
rect 30380 8910 30432 8916
rect 30286 8664 30342 8673
rect 30286 8599 30342 8608
rect 30196 8560 30248 8566
rect 30196 8502 30248 8508
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 30012 8356 30064 8362
rect 30012 8298 30064 8304
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 30024 8106 30052 8298
rect 30208 8276 30236 8502
rect 30288 8424 30340 8430
rect 30286 8392 30288 8401
rect 30340 8392 30342 8401
rect 30286 8327 30342 8336
rect 30208 8248 30328 8276
rect 29932 8078 30052 8106
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 29840 7750 29868 7822
rect 29828 7744 29880 7750
rect 29828 7686 29880 7692
rect 29828 6860 29880 6866
rect 29828 6802 29880 6808
rect 29840 6497 29868 6802
rect 29932 6662 29960 8078
rect 30010 7984 30066 7993
rect 30010 7919 30066 7928
rect 29920 6656 29972 6662
rect 29920 6598 29972 6604
rect 29826 6488 29882 6497
rect 29826 6423 29882 6432
rect 29828 6384 29880 6390
rect 29828 6326 29880 6332
rect 29840 4622 29868 6326
rect 29918 5672 29974 5681
rect 29918 5607 29974 5616
rect 29828 4616 29880 4622
rect 29828 4558 29880 4564
rect 29840 4214 29868 4558
rect 29828 4208 29880 4214
rect 29828 4150 29880 4156
rect 29736 3732 29788 3738
rect 29736 3674 29788 3680
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 29196 2650 29224 2994
rect 29184 2644 29236 2650
rect 29184 2586 29236 2592
rect 29932 2446 29960 5607
rect 30024 4826 30052 7919
rect 30300 7818 30328 8248
rect 30288 7812 30340 7818
rect 30288 7754 30340 7760
rect 30102 7440 30158 7449
rect 30102 7375 30158 7384
rect 30116 7274 30144 7375
rect 30300 7342 30328 7754
rect 30288 7336 30340 7342
rect 30288 7278 30340 7284
rect 30104 7268 30156 7274
rect 30104 7210 30156 7216
rect 30196 7268 30248 7274
rect 30196 7210 30248 7216
rect 30208 6866 30236 7210
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 30392 6730 30420 8910
rect 30484 8566 30512 13926
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30576 11150 30604 11630
rect 30668 11354 30696 17138
rect 30944 16794 30972 17190
rect 31024 17138 31076 17144
rect 31576 17128 31628 17134
rect 31576 17070 31628 17076
rect 31588 16794 31616 17070
rect 30932 16788 30984 16794
rect 30932 16730 30984 16736
rect 31576 16788 31628 16794
rect 31576 16730 31628 16736
rect 31588 16697 31616 16730
rect 31574 16688 31630 16697
rect 31574 16623 31630 16632
rect 31208 16584 31260 16590
rect 31208 16526 31260 16532
rect 31220 16182 31248 16526
rect 31300 16448 31352 16454
rect 31300 16390 31352 16396
rect 31208 16176 31260 16182
rect 31208 16118 31260 16124
rect 31024 16108 31076 16114
rect 31024 16050 31076 16056
rect 30840 15700 30892 15706
rect 30840 15642 30892 15648
rect 30852 15502 30880 15642
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 31036 15434 31064 16050
rect 31116 15972 31168 15978
rect 31116 15914 31168 15920
rect 30932 15428 30984 15434
rect 30932 15370 30984 15376
rect 31024 15428 31076 15434
rect 31024 15370 31076 15376
rect 30944 15026 30972 15370
rect 31128 15094 31156 15914
rect 31220 15706 31248 16118
rect 31312 16114 31340 16390
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31208 15700 31260 15706
rect 31208 15642 31260 15648
rect 31312 15366 31340 16050
rect 31404 15502 31432 16050
rect 31392 15496 31444 15502
rect 31392 15438 31444 15444
rect 31300 15360 31352 15366
rect 31300 15302 31352 15308
rect 31116 15088 31168 15094
rect 31116 15030 31168 15036
rect 31392 15088 31444 15094
rect 31392 15030 31444 15036
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 31404 14414 31432 15030
rect 31852 15020 31904 15026
rect 31852 14962 31904 14968
rect 31760 14816 31812 14822
rect 31760 14758 31812 14764
rect 31116 14408 31168 14414
rect 31116 14350 31168 14356
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31576 14408 31628 14414
rect 31576 14350 31628 14356
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 31036 13841 31064 13874
rect 31022 13832 31078 13841
rect 31022 13767 31078 13776
rect 31128 13734 31156 14350
rect 31300 14068 31352 14074
rect 31300 14010 31352 14016
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31312 13530 31340 14010
rect 31300 13524 31352 13530
rect 31300 13466 31352 13472
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30748 13252 30800 13258
rect 30748 13194 30800 13200
rect 30760 12646 30788 13194
rect 30748 12640 30800 12646
rect 30748 12582 30800 12588
rect 30760 12238 30788 12582
rect 30748 12232 30800 12238
rect 30748 12174 30800 12180
rect 30748 12096 30800 12102
rect 30748 12038 30800 12044
rect 30760 11762 30788 12038
rect 30748 11756 30800 11762
rect 30748 11698 30800 11704
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30576 10266 30604 11086
rect 30748 10804 30800 10810
rect 30748 10746 30800 10752
rect 30564 10260 30616 10266
rect 30564 10202 30616 10208
rect 30564 10056 30616 10062
rect 30564 9998 30616 10004
rect 30576 9518 30604 9998
rect 30564 9512 30616 9518
rect 30564 9454 30616 9460
rect 30656 9444 30708 9450
rect 30656 9386 30708 9392
rect 30472 8560 30524 8566
rect 30472 8502 30524 8508
rect 30472 8424 30524 8430
rect 30524 8384 30604 8412
rect 30472 8366 30524 8372
rect 30472 7744 30524 7750
rect 30472 7686 30524 7692
rect 30484 7410 30512 7686
rect 30472 7404 30524 7410
rect 30472 7346 30524 7352
rect 30576 6798 30604 8384
rect 30668 7750 30696 9386
rect 30656 7744 30708 7750
rect 30656 7686 30708 7692
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30380 6724 30432 6730
rect 30380 6666 30432 6672
rect 30392 6254 30420 6666
rect 30576 6322 30604 6734
rect 30760 6390 30788 10746
rect 30852 9178 30880 13262
rect 31024 12640 31076 12646
rect 31024 12582 31076 12588
rect 31036 11830 31064 12582
rect 31588 12434 31616 14350
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31680 13462 31708 13874
rect 31772 13870 31800 14758
rect 31760 13864 31812 13870
rect 31760 13806 31812 13812
rect 31668 13456 31720 13462
rect 31668 13398 31720 13404
rect 31496 12406 31616 12434
rect 31024 11824 31076 11830
rect 31024 11766 31076 11772
rect 31036 11665 31064 11766
rect 31022 11656 31078 11665
rect 31022 11591 31078 11600
rect 31116 11620 31168 11626
rect 31300 11620 31352 11626
rect 31168 11580 31300 11608
rect 31116 11562 31168 11568
rect 31300 11562 31352 11568
rect 30932 11144 30984 11150
rect 31208 11144 31260 11150
rect 30932 11086 30984 11092
rect 31128 11104 31208 11132
rect 30944 10810 30972 11086
rect 30932 10804 30984 10810
rect 30932 10746 30984 10752
rect 30930 10568 30986 10577
rect 30930 10503 30986 10512
rect 30944 10470 30972 10503
rect 30932 10464 30984 10470
rect 30932 10406 30984 10412
rect 30930 10160 30986 10169
rect 30930 10095 30986 10104
rect 30944 9674 30972 10095
rect 30944 9646 31064 9674
rect 31128 9654 31156 11104
rect 31208 11086 31260 11092
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 31208 11008 31260 11014
rect 31208 10950 31260 10956
rect 31220 10470 31248 10950
rect 31300 10804 31352 10810
rect 31300 10746 31352 10752
rect 31208 10464 31260 10470
rect 31208 10406 31260 10412
rect 31312 10062 31340 10746
rect 31300 10056 31352 10062
rect 31206 10024 31262 10033
rect 31300 9998 31352 10004
rect 31206 9959 31208 9968
rect 31260 9959 31262 9968
rect 31208 9930 31260 9936
rect 31300 9920 31352 9926
rect 31300 9862 31352 9868
rect 30932 9580 30984 9586
rect 30932 9522 30984 9528
rect 30840 9172 30892 9178
rect 30840 9114 30892 9120
rect 30840 8832 30892 8838
rect 30944 8809 30972 9522
rect 30840 8774 30892 8780
rect 30930 8800 30986 8809
rect 30852 8430 30880 8774
rect 30930 8735 30986 8744
rect 30840 8424 30892 8430
rect 30840 8366 30892 8372
rect 30840 7268 30892 7274
rect 30840 7210 30892 7216
rect 30852 7002 30880 7210
rect 30840 6996 30892 7002
rect 30840 6938 30892 6944
rect 30944 6458 30972 8735
rect 31036 6798 31064 9646
rect 31116 9648 31168 9654
rect 31116 9590 31168 9596
rect 31208 9580 31260 9586
rect 31208 9522 31260 9528
rect 31116 9444 31168 9450
rect 31116 9386 31168 9392
rect 31128 7750 31156 9386
rect 31116 7744 31168 7750
rect 31116 7686 31168 7692
rect 31128 7449 31156 7686
rect 31220 7585 31248 9522
rect 31312 9382 31340 9862
rect 31300 9376 31352 9382
rect 31300 9318 31352 9324
rect 31404 8974 31432 11018
rect 31496 9160 31524 12406
rect 31574 11656 31630 11665
rect 31574 11591 31630 11600
rect 31588 9654 31616 11591
rect 31680 11558 31708 13398
rect 31864 12986 31892 14962
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 31852 12164 31904 12170
rect 31852 12106 31904 12112
rect 31864 11830 31892 12106
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 31852 11824 31904 11830
rect 31852 11766 31904 11772
rect 31668 11552 31720 11558
rect 31668 11494 31720 11500
rect 31680 11218 31708 11494
rect 31850 11248 31906 11257
rect 31668 11212 31720 11218
rect 31850 11183 31906 11192
rect 31668 11154 31720 11160
rect 31668 11008 31720 11014
rect 31864 10996 31892 11183
rect 31956 11121 31984 12038
rect 32048 11234 32076 57326
rect 43732 57254 43760 57394
rect 43720 57248 43772 57254
rect 43720 57190 43772 57196
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 40408 56840 40460 56846
rect 40408 56782 40460 56788
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 40040 26512 40092 26518
rect 40040 26454 40092 26460
rect 38476 26308 38528 26314
rect 38476 26250 38528 26256
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 37740 25288 37792 25294
rect 37740 25230 37792 25236
rect 38016 25288 38068 25294
rect 38016 25230 38068 25236
rect 38200 25288 38252 25294
rect 38200 25230 38252 25236
rect 37188 25220 37240 25226
rect 37188 25162 37240 25168
rect 37200 24954 37228 25162
rect 37464 25152 37516 25158
rect 37464 25094 37516 25100
rect 37188 24948 37240 24954
rect 37188 24890 37240 24896
rect 37476 24886 37504 25094
rect 37464 24880 37516 24886
rect 37464 24822 37516 24828
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 36452 24812 36504 24818
rect 36452 24754 36504 24760
rect 34796 24744 34848 24750
rect 34796 24686 34848 24692
rect 34808 24274 34836 24686
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 24268 34848 24274
rect 34796 24210 34848 24216
rect 32496 24200 32548 24206
rect 32496 24142 32548 24148
rect 35256 24200 35308 24206
rect 35360 24188 35388 24754
rect 36360 24744 36412 24750
rect 36360 24686 36412 24692
rect 35624 24676 35676 24682
rect 35624 24618 35676 24624
rect 35636 24410 35664 24618
rect 35624 24404 35676 24410
rect 35624 24346 35676 24352
rect 36268 24404 36320 24410
rect 36268 24346 36320 24352
rect 35308 24160 35388 24188
rect 35256 24142 35308 24148
rect 32508 23186 32536 24142
rect 35268 23866 35296 24142
rect 35256 23860 35308 23866
rect 35256 23802 35308 23808
rect 34520 23656 34572 23662
rect 34520 23598 34572 23604
rect 34532 23322 34560 23598
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34520 23316 34572 23322
rect 34520 23258 34572 23264
rect 32496 23180 32548 23186
rect 32496 23122 32548 23128
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 32140 22030 32168 23054
rect 34704 23044 34756 23050
rect 34704 22986 34756 22992
rect 33968 22976 34020 22982
rect 33968 22918 34020 22924
rect 33980 22642 34008 22918
rect 33968 22636 34020 22642
rect 33968 22578 34020 22584
rect 32588 22160 32640 22166
rect 32588 22102 32640 22108
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 32140 21690 32168 21966
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 32220 21548 32272 21554
rect 32220 21490 32272 21496
rect 32232 20806 32260 21490
rect 32600 21486 32628 22102
rect 34520 22092 34572 22098
rect 34520 22034 34572 22040
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 32588 21480 32640 21486
rect 32588 21422 32640 21428
rect 32956 21480 33008 21486
rect 32956 21422 33008 21428
rect 32312 21412 32364 21418
rect 32312 21354 32364 21360
rect 32324 21146 32352 21354
rect 32968 21350 32996 21422
rect 32956 21344 33008 21350
rect 32956 21286 33008 21292
rect 32312 21140 32364 21146
rect 32312 21082 32364 21088
rect 32968 20874 32996 21286
rect 33336 21146 33364 21966
rect 33692 21548 33744 21554
rect 33692 21490 33744 21496
rect 33324 21140 33376 21146
rect 33324 21082 33376 21088
rect 33704 21078 33732 21490
rect 33784 21344 33836 21350
rect 33784 21286 33836 21292
rect 33692 21072 33744 21078
rect 33692 21014 33744 21020
rect 32956 20868 33008 20874
rect 32956 20810 33008 20816
rect 33508 20868 33560 20874
rect 33508 20810 33560 20816
rect 32220 20800 32272 20806
rect 32220 20742 32272 20748
rect 32232 20398 32260 20742
rect 33232 20460 33284 20466
rect 33232 20402 33284 20408
rect 33416 20460 33468 20466
rect 33416 20402 33468 20408
rect 32220 20392 32272 20398
rect 32220 20334 32272 20340
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32232 19378 32260 19790
rect 33244 19786 33272 20402
rect 33428 19922 33456 20402
rect 33520 20058 33548 20810
rect 33704 20602 33732 21014
rect 33796 21010 33824 21286
rect 33784 21004 33836 21010
rect 33784 20946 33836 20952
rect 34532 20942 34560 22034
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 34532 20602 34560 20878
rect 33692 20596 33744 20602
rect 33692 20538 33744 20544
rect 34520 20596 34572 20602
rect 34520 20538 34572 20544
rect 33784 20460 33836 20466
rect 33784 20402 33836 20408
rect 33508 20052 33560 20058
rect 33508 19994 33560 20000
rect 33416 19916 33468 19922
rect 33416 19858 33468 19864
rect 33796 19786 33824 20402
rect 34612 19848 34664 19854
rect 34612 19790 34664 19796
rect 33232 19780 33284 19786
rect 33232 19722 33284 19728
rect 33784 19780 33836 19786
rect 33784 19722 33836 19728
rect 32680 19712 32732 19718
rect 32680 19654 32732 19660
rect 32692 19446 32720 19654
rect 32680 19440 32732 19446
rect 32680 19382 32732 19388
rect 32220 19372 32272 19378
rect 32220 19314 32272 19320
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 32232 18766 32260 19314
rect 32128 18760 32180 18766
rect 32128 18702 32180 18708
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32140 17610 32168 18702
rect 32220 18216 32272 18222
rect 32220 18158 32272 18164
rect 32128 17604 32180 17610
rect 32128 17546 32180 17552
rect 32232 15502 32260 18158
rect 32312 17740 32364 17746
rect 32312 17682 32364 17688
rect 32324 17134 32352 17682
rect 32416 17678 32444 19314
rect 32496 19304 32548 19310
rect 32496 19246 32548 19252
rect 32508 18970 32536 19246
rect 32496 18964 32548 18970
rect 32496 18906 32548 18912
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 32692 17678 32720 18702
rect 33152 18290 33180 19314
rect 33244 19310 33272 19722
rect 33232 19304 33284 19310
rect 33232 19246 33284 19252
rect 33232 18828 33284 18834
rect 33232 18770 33284 18776
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32956 18284 33008 18290
rect 32956 18226 33008 18232
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 32404 17672 32456 17678
rect 32404 17614 32456 17620
rect 32680 17672 32732 17678
rect 32680 17614 32732 17620
rect 32312 17128 32364 17134
rect 32312 17070 32364 17076
rect 32324 16726 32352 17070
rect 32312 16720 32364 16726
rect 32312 16662 32364 16668
rect 32220 15496 32272 15502
rect 32220 15438 32272 15444
rect 32232 15026 32260 15438
rect 32312 15428 32364 15434
rect 32312 15370 32364 15376
rect 32220 15020 32272 15026
rect 32220 14962 32272 14968
rect 32324 14958 32352 15370
rect 32312 14952 32364 14958
rect 32312 14894 32364 14900
rect 32324 14618 32352 14894
rect 32416 14618 32444 17614
rect 32496 15972 32548 15978
rect 32496 15914 32548 15920
rect 32508 14890 32536 15914
rect 32692 15586 32720 17614
rect 32784 16454 32812 18226
rect 32968 17134 32996 18226
rect 33152 17338 33180 18226
rect 33244 17882 33272 18770
rect 33796 17882 33824 19722
rect 34624 19514 34652 19790
rect 34716 19514 34744 22986
rect 34796 22636 34848 22642
rect 34796 22578 34848 22584
rect 34808 22234 34836 22578
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 22228 34848 22234
rect 34796 22170 34848 22176
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34612 19508 34664 19514
rect 34532 19446 34560 19477
rect 34612 19450 34664 19456
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34520 19440 34572 19446
rect 34572 19388 34928 19394
rect 34520 19382 34928 19388
rect 34532 19378 34928 19382
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34532 19372 34940 19378
rect 34532 19366 34888 19372
rect 33232 17876 33284 17882
rect 33232 17818 33284 17824
rect 33784 17876 33836 17882
rect 33784 17818 33836 17824
rect 33244 17678 33272 17818
rect 34060 17740 34112 17746
rect 34060 17682 34112 17688
rect 33232 17672 33284 17678
rect 33232 17614 33284 17620
rect 33692 17672 33744 17678
rect 33692 17614 33744 17620
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 32956 17128 33008 17134
rect 32956 17070 33008 17076
rect 33140 16652 33192 16658
rect 33140 16594 33192 16600
rect 33048 16584 33100 16590
rect 33048 16526 33100 16532
rect 32956 16516 33008 16522
rect 32956 16458 33008 16464
rect 32772 16448 32824 16454
rect 32772 16390 32824 16396
rect 32772 16040 32824 16046
rect 32772 15982 32824 15988
rect 32784 15706 32812 15982
rect 32772 15700 32824 15706
rect 32772 15642 32824 15648
rect 32692 15558 32812 15586
rect 32680 14952 32732 14958
rect 32680 14894 32732 14900
rect 32496 14884 32548 14890
rect 32496 14826 32548 14832
rect 32588 14884 32640 14890
rect 32588 14826 32640 14832
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32404 14612 32456 14618
rect 32404 14554 32456 14560
rect 32600 14414 32628 14826
rect 32692 14550 32720 14894
rect 32680 14544 32732 14550
rect 32680 14486 32732 14492
rect 32312 14408 32364 14414
rect 32312 14350 32364 14356
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 32588 14408 32640 14414
rect 32784 14396 32812 15558
rect 32968 15502 32996 16458
rect 33060 16454 33088 16526
rect 33048 16448 33100 16454
rect 33048 16390 33100 16396
rect 33060 16250 33088 16390
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 32956 15496 33008 15502
rect 32956 15438 33008 15444
rect 32864 14816 32916 14822
rect 32864 14758 32916 14764
rect 32876 14414 32904 14758
rect 32588 14350 32640 14356
rect 32692 14368 32812 14396
rect 32864 14408 32916 14414
rect 32220 13864 32272 13870
rect 32220 13806 32272 13812
rect 32128 13728 32180 13734
rect 32128 13670 32180 13676
rect 32140 13530 32168 13670
rect 32128 13524 32180 13530
rect 32128 13466 32180 13472
rect 32048 11206 32168 11234
rect 32036 11144 32088 11150
rect 31942 11112 31998 11121
rect 32036 11086 32088 11092
rect 31942 11047 31998 11056
rect 31864 10968 31984 10996
rect 31668 10950 31720 10956
rect 31680 10062 31708 10950
rect 31956 10690 31984 10968
rect 32048 10810 32076 11086
rect 32036 10804 32088 10810
rect 32036 10746 32088 10752
rect 31760 10668 31812 10674
rect 31956 10662 32076 10690
rect 31760 10610 31812 10616
rect 31772 10266 31800 10610
rect 31760 10260 31812 10266
rect 31760 10202 31812 10208
rect 31758 10160 31814 10169
rect 31758 10095 31814 10104
rect 31668 10056 31720 10062
rect 31668 9998 31720 10004
rect 31680 9926 31708 9998
rect 31668 9920 31720 9926
rect 31668 9862 31720 9868
rect 31576 9648 31628 9654
rect 31576 9590 31628 9596
rect 31576 9172 31628 9178
rect 31496 9132 31576 9160
rect 31392 8968 31444 8974
rect 31392 8910 31444 8916
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 31206 7576 31262 7585
rect 31206 7511 31262 7520
rect 31114 7440 31170 7449
rect 31114 7375 31170 7384
rect 31116 6928 31168 6934
rect 31116 6870 31168 6876
rect 31128 6798 31156 6870
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 30932 6452 30984 6458
rect 30932 6394 30984 6400
rect 30748 6384 30800 6390
rect 30748 6326 30800 6332
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30380 6248 30432 6254
rect 30380 6190 30432 6196
rect 30576 5710 30604 6258
rect 30760 5846 30788 6326
rect 30748 5840 30800 5846
rect 30748 5782 30800 5788
rect 30196 5704 30248 5710
rect 30196 5646 30248 5652
rect 30564 5704 30616 5710
rect 30564 5646 30616 5652
rect 30102 5400 30158 5409
rect 30102 5335 30104 5344
rect 30156 5335 30158 5344
rect 30104 5306 30156 5312
rect 30208 5302 30236 5646
rect 30196 5296 30248 5302
rect 30196 5238 30248 5244
rect 30760 5234 30788 5782
rect 30748 5228 30800 5234
rect 30748 5170 30800 5176
rect 30472 5092 30524 5098
rect 30472 5034 30524 5040
rect 30196 5024 30248 5030
rect 30196 4966 30248 4972
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 30024 3738 30052 4762
rect 30208 4690 30236 4966
rect 30196 4684 30248 4690
rect 30196 4626 30248 4632
rect 30208 4264 30236 4626
rect 30208 4236 30328 4264
rect 30300 4146 30328 4236
rect 30196 4140 30248 4146
rect 30196 4082 30248 4088
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 30208 3534 30236 4082
rect 30300 3942 30328 4082
rect 30288 3936 30340 3942
rect 30288 3878 30340 3884
rect 30300 3602 30328 3878
rect 30288 3596 30340 3602
rect 30288 3538 30340 3544
rect 30196 3528 30248 3534
rect 30196 3470 30248 3476
rect 30208 3126 30236 3470
rect 30196 3120 30248 3126
rect 30196 3062 30248 3068
rect 30300 2854 30328 3538
rect 30484 2922 30512 5034
rect 31128 4826 31156 6734
rect 31116 4820 31168 4826
rect 31116 4762 31168 4768
rect 31220 4758 31248 7511
rect 31312 7410 31340 8570
rect 31404 8537 31432 8774
rect 31390 8528 31446 8537
rect 31390 8463 31392 8472
rect 31444 8463 31446 8472
rect 31392 8434 31444 8440
rect 31300 7404 31352 7410
rect 31300 7346 31352 7352
rect 31404 6866 31432 8434
rect 31496 7886 31524 9132
rect 31576 9114 31628 9120
rect 31576 9036 31628 9042
rect 31576 8978 31628 8984
rect 31484 7880 31536 7886
rect 31484 7822 31536 7828
rect 31496 7410 31524 7822
rect 31588 7546 31616 8978
rect 31680 8838 31708 9862
rect 31772 9110 31800 10095
rect 31944 9988 31996 9994
rect 31944 9930 31996 9936
rect 31760 9104 31812 9110
rect 31760 9046 31812 9052
rect 31668 8832 31720 8838
rect 31668 8774 31720 8780
rect 31852 8832 31904 8838
rect 31852 8774 31904 8780
rect 31864 8498 31892 8774
rect 31852 8492 31904 8498
rect 31852 8434 31904 8440
rect 31758 7984 31814 7993
rect 31758 7919 31814 7928
rect 31772 7886 31800 7919
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31576 7540 31628 7546
rect 31576 7482 31628 7488
rect 31666 7440 31722 7449
rect 31484 7404 31536 7410
rect 31666 7375 31722 7384
rect 31484 7346 31536 7352
rect 31392 6860 31444 6866
rect 31392 6802 31444 6808
rect 31496 6390 31524 7346
rect 31680 7206 31708 7375
rect 31668 7200 31720 7206
rect 31668 7142 31720 7148
rect 31864 7041 31892 8434
rect 31666 7032 31722 7041
rect 31666 6967 31722 6976
rect 31850 7032 31906 7041
rect 31850 6967 31906 6976
rect 31680 6662 31708 6967
rect 31852 6792 31904 6798
rect 31956 6780 31984 9930
rect 32048 9518 32076 10662
rect 32140 9625 32168 11206
rect 32232 10538 32260 13806
rect 32324 11354 32352 14350
rect 32508 14074 32536 14350
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 32600 12782 32628 13874
rect 32496 12776 32548 12782
rect 32496 12718 32548 12724
rect 32588 12776 32640 12782
rect 32588 12718 32640 12724
rect 32508 12442 32536 12718
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 32404 12368 32456 12374
rect 32404 12310 32456 12316
rect 32416 12102 32444 12310
rect 32404 12096 32456 12102
rect 32404 12038 32456 12044
rect 32312 11348 32364 11354
rect 32312 11290 32364 11296
rect 32310 11112 32366 11121
rect 32310 11047 32366 11056
rect 32220 10532 32272 10538
rect 32220 10474 32272 10480
rect 32324 10418 32352 11047
rect 32232 10390 32352 10418
rect 32232 10062 32260 10390
rect 32416 10282 32444 12038
rect 32494 11792 32550 11801
rect 32494 11727 32496 11736
rect 32548 11727 32550 11736
rect 32496 11698 32548 11704
rect 32496 11620 32548 11626
rect 32496 11562 32548 11568
rect 32324 10254 32444 10282
rect 32220 10056 32272 10062
rect 32220 9998 32272 10004
rect 32126 9616 32182 9625
rect 32126 9551 32182 9560
rect 32036 9512 32088 9518
rect 32036 9454 32088 9460
rect 32048 8906 32076 9454
rect 32232 8922 32260 9998
rect 32324 9489 32352 10254
rect 32404 9648 32456 9654
rect 32404 9590 32456 9596
rect 32310 9480 32366 9489
rect 32310 9415 32366 9424
rect 32036 8900 32088 8906
rect 32036 8842 32088 8848
rect 32140 8894 32260 8922
rect 32310 8936 32366 8945
rect 32140 8537 32168 8894
rect 32310 8871 32312 8880
rect 32364 8871 32366 8880
rect 32312 8842 32364 8848
rect 32220 8832 32272 8838
rect 32220 8774 32272 8780
rect 32126 8528 32182 8537
rect 32126 8463 32182 8472
rect 32034 8256 32090 8265
rect 32034 8191 32090 8200
rect 32048 7410 32076 8191
rect 32140 7886 32168 8463
rect 32128 7880 32180 7886
rect 32128 7822 32180 7828
rect 32036 7404 32088 7410
rect 32036 7346 32088 7352
rect 31904 6752 31984 6780
rect 31852 6734 31904 6740
rect 31668 6656 31720 6662
rect 31668 6598 31720 6604
rect 31484 6384 31536 6390
rect 31484 6326 31536 6332
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31392 6316 31444 6322
rect 31392 6258 31444 6264
rect 31312 5234 31340 6258
rect 31404 6089 31432 6258
rect 31390 6080 31446 6089
rect 31390 6015 31446 6024
rect 31390 5944 31446 5953
rect 31390 5879 31392 5888
rect 31444 5879 31446 5888
rect 31392 5850 31444 5856
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 31864 5370 31892 5646
rect 31852 5364 31904 5370
rect 31852 5306 31904 5312
rect 31300 5228 31352 5234
rect 31300 5170 31352 5176
rect 31484 5228 31536 5234
rect 31484 5170 31536 5176
rect 31852 5228 31904 5234
rect 31956 5216 31984 6752
rect 32128 6792 32180 6798
rect 32128 6734 32180 6740
rect 32140 6497 32168 6734
rect 32126 6488 32182 6497
rect 32126 6423 32128 6432
rect 32180 6423 32182 6432
rect 32128 6394 32180 6400
rect 32140 6363 32168 6394
rect 32232 5914 32260 8774
rect 32324 7818 32352 8842
rect 32312 7812 32364 7818
rect 32312 7754 32364 7760
rect 32220 5908 32272 5914
rect 32220 5850 32272 5856
rect 32036 5772 32088 5778
rect 32036 5714 32088 5720
rect 31904 5188 31984 5216
rect 31852 5170 31904 5176
rect 31208 4752 31260 4758
rect 31208 4694 31260 4700
rect 31208 4548 31260 4554
rect 31208 4490 31260 4496
rect 31220 3398 31248 4490
rect 31312 3738 31340 5170
rect 31496 4622 31524 5170
rect 31852 4752 31904 4758
rect 31852 4694 31904 4700
rect 31484 4616 31536 4622
rect 31484 4558 31536 4564
rect 31864 4282 31892 4694
rect 31852 4276 31904 4282
rect 31852 4218 31904 4224
rect 31484 4140 31536 4146
rect 31484 4082 31536 4088
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 31208 3392 31260 3398
rect 31208 3334 31260 3340
rect 31220 3126 31248 3334
rect 31496 3126 31524 4082
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 31864 3738 31892 3878
rect 31852 3732 31904 3738
rect 31852 3674 31904 3680
rect 31208 3120 31260 3126
rect 31208 3062 31260 3068
rect 31484 3120 31536 3126
rect 31484 3062 31536 3068
rect 31220 2922 31248 3062
rect 32048 3058 32076 5714
rect 32324 5302 32352 7754
rect 32312 5296 32364 5302
rect 32312 5238 32364 5244
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 32324 4622 32352 4966
rect 32312 4616 32364 4622
rect 32312 4558 32364 4564
rect 32220 4072 32272 4078
rect 32220 4014 32272 4020
rect 32232 3738 32260 4014
rect 32220 3732 32272 3738
rect 32220 3674 32272 3680
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 30472 2916 30524 2922
rect 30472 2858 30524 2864
rect 31208 2916 31260 2922
rect 31208 2858 31260 2864
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 31024 2848 31076 2854
rect 31024 2790 31076 2796
rect 31036 2650 31064 2790
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 31220 2446 31248 2858
rect 32324 2854 32352 4558
rect 32416 4214 32444 9590
rect 32508 8945 32536 11562
rect 32588 10532 32640 10538
rect 32588 10474 32640 10480
rect 32494 8936 32550 8945
rect 32494 8871 32550 8880
rect 32508 8566 32536 8871
rect 32496 8560 32548 8566
rect 32496 8502 32548 8508
rect 32496 7880 32548 7886
rect 32496 7822 32548 7828
rect 32508 7546 32536 7822
rect 32496 7540 32548 7546
rect 32496 7482 32548 7488
rect 32494 7440 32550 7449
rect 32494 7375 32550 7384
rect 32508 7342 32536 7375
rect 32496 7336 32548 7342
rect 32496 7278 32548 7284
rect 32494 6760 32550 6769
rect 32494 6695 32550 6704
rect 32508 6662 32536 6695
rect 32496 6656 32548 6662
rect 32496 6598 32548 6604
rect 32600 6458 32628 10474
rect 32692 9654 32720 14368
rect 32864 14350 32916 14356
rect 32956 13932 33008 13938
rect 32956 13874 33008 13880
rect 32864 12708 32916 12714
rect 32864 12650 32916 12656
rect 32770 11112 32826 11121
rect 32770 11047 32772 11056
rect 32824 11047 32826 11056
rect 32772 11018 32824 11024
rect 32784 10742 32812 11018
rect 32772 10736 32824 10742
rect 32772 10678 32824 10684
rect 32772 10600 32824 10606
rect 32772 10542 32824 10548
rect 32784 10130 32812 10542
rect 32772 10124 32824 10130
rect 32772 10066 32824 10072
rect 32772 9920 32824 9926
rect 32772 9862 32824 9868
rect 32680 9648 32732 9654
rect 32680 9590 32732 9596
rect 32784 8809 32812 9862
rect 32876 9178 32904 12650
rect 32968 11354 32996 13874
rect 33048 13388 33100 13394
rect 33048 13330 33100 13336
rect 33060 12238 33088 13330
rect 33152 12442 33180 16594
rect 33704 16250 33732 17614
rect 34072 17338 34100 17682
rect 34060 17332 34112 17338
rect 34060 17274 34112 17280
rect 33784 17196 33836 17202
rect 33784 17138 33836 17144
rect 34152 17196 34204 17202
rect 34152 17138 34204 17144
rect 33796 16590 33824 17138
rect 34164 16590 34192 17138
rect 33784 16584 33836 16590
rect 33784 16526 33836 16532
rect 34152 16584 34204 16590
rect 34152 16526 34204 16532
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33416 16108 33468 16114
rect 33416 16050 33468 16056
rect 33324 16040 33376 16046
rect 33324 15982 33376 15988
rect 33336 15502 33364 15982
rect 33324 15496 33376 15502
rect 33324 15438 33376 15444
rect 33336 13870 33364 15438
rect 33428 15366 33456 16050
rect 34164 15502 34192 16526
rect 34440 16250 34468 19314
rect 34532 18834 34560 19366
rect 34888 19314 34940 19320
rect 34796 19304 34848 19310
rect 34796 19246 34848 19252
rect 34808 18970 34836 19246
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34796 18964 34848 18970
rect 34796 18906 34848 18912
rect 34520 18828 34572 18834
rect 34520 18770 34572 18776
rect 34532 17814 34560 18770
rect 35360 18426 35388 23054
rect 35532 22024 35584 22030
rect 35532 21966 35584 21972
rect 35440 21956 35492 21962
rect 35440 21898 35492 21904
rect 35452 21622 35480 21898
rect 35440 21616 35492 21622
rect 35440 21558 35492 21564
rect 35544 21554 35572 21966
rect 35532 21548 35584 21554
rect 35532 21490 35584 21496
rect 35544 21078 35572 21490
rect 35532 21072 35584 21078
rect 35532 21014 35584 21020
rect 35532 20936 35584 20942
rect 35636 20924 35664 24346
rect 35900 23724 35952 23730
rect 35900 23666 35952 23672
rect 35912 23322 35940 23666
rect 35900 23316 35952 23322
rect 35900 23258 35952 23264
rect 36280 23118 36308 24346
rect 36372 23866 36400 24686
rect 36464 24206 36492 24754
rect 37476 24410 37504 24822
rect 37752 24614 37780 25230
rect 37740 24608 37792 24614
rect 37740 24550 37792 24556
rect 37464 24404 37516 24410
rect 37464 24346 37516 24352
rect 36452 24200 36504 24206
rect 36452 24142 36504 24148
rect 36360 23860 36412 23866
rect 36360 23802 36412 23808
rect 36464 23798 36492 24142
rect 36452 23792 36504 23798
rect 36452 23734 36504 23740
rect 36464 23186 36492 23734
rect 36452 23180 36504 23186
rect 36452 23122 36504 23128
rect 37464 23180 37516 23186
rect 37464 23122 37516 23128
rect 36268 23112 36320 23118
rect 36268 23054 36320 23060
rect 35900 21548 35952 21554
rect 35900 21490 35952 21496
rect 35912 21146 35940 21490
rect 35900 21140 35952 21146
rect 35900 21082 35952 21088
rect 35716 21004 35768 21010
rect 35716 20946 35768 20952
rect 35584 20896 35664 20924
rect 35532 20878 35584 20884
rect 35440 20460 35492 20466
rect 35440 20402 35492 20408
rect 35452 20058 35480 20402
rect 35440 20052 35492 20058
rect 35440 19994 35492 20000
rect 35544 19938 35572 20878
rect 35624 20800 35676 20806
rect 35624 20742 35676 20748
rect 35452 19910 35572 19938
rect 35256 18420 35308 18426
rect 35256 18362 35308 18368
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35268 18086 35296 18362
rect 35256 18080 35308 18086
rect 35256 18022 35308 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35452 17882 35480 19910
rect 35532 19372 35584 19378
rect 35532 19314 35584 19320
rect 35440 17876 35492 17882
rect 35440 17818 35492 17824
rect 34520 17808 34572 17814
rect 34520 17750 34572 17756
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34532 16454 34560 17614
rect 35544 17338 35572 19314
rect 35636 18970 35664 20742
rect 35624 18964 35676 18970
rect 35624 18906 35676 18912
rect 35624 18692 35676 18698
rect 35624 18634 35676 18640
rect 35636 17338 35664 18634
rect 35532 17332 35584 17338
rect 35532 17274 35584 17280
rect 35624 17332 35676 17338
rect 35624 17274 35676 17280
rect 34704 17196 34756 17202
rect 34704 17138 34756 17144
rect 34612 17128 34664 17134
rect 34612 17070 34664 17076
rect 34520 16448 34572 16454
rect 34520 16390 34572 16396
rect 34428 16244 34480 16250
rect 34428 16186 34480 16192
rect 34152 15496 34204 15502
rect 34152 15438 34204 15444
rect 33416 15360 33468 15366
rect 33416 15302 33468 15308
rect 34336 15360 34388 15366
rect 34336 15302 34388 15308
rect 33428 14618 33456 15302
rect 34348 15026 34376 15302
rect 34428 15088 34480 15094
rect 34428 15030 34480 15036
rect 34336 15020 34388 15026
rect 34336 14962 34388 14968
rect 33416 14612 33468 14618
rect 33416 14554 33468 14560
rect 33784 14476 33836 14482
rect 33704 14436 33784 14464
rect 33600 14340 33652 14346
rect 33600 14282 33652 14288
rect 33612 14074 33640 14282
rect 33704 14074 33732 14436
rect 33784 14418 33836 14424
rect 33876 14272 33928 14278
rect 33876 14214 33928 14220
rect 33968 14272 34020 14278
rect 33968 14214 34020 14220
rect 33600 14068 33652 14074
rect 33600 14010 33652 14016
rect 33692 14068 33744 14074
rect 33692 14010 33744 14016
rect 33416 13932 33468 13938
rect 33416 13874 33468 13880
rect 33324 13864 33376 13870
rect 33324 13806 33376 13812
rect 33232 13320 33284 13326
rect 33232 13262 33284 13268
rect 33140 12436 33192 12442
rect 33140 12378 33192 12384
rect 33048 12232 33100 12238
rect 33048 12174 33100 12180
rect 33060 11762 33088 12174
rect 33048 11756 33100 11762
rect 33048 11698 33100 11704
rect 33244 11642 33272 13262
rect 33428 12986 33456 13874
rect 33508 13796 33560 13802
rect 33508 13738 33560 13744
rect 33520 13190 33548 13738
rect 33600 13456 33652 13462
rect 33600 13398 33652 13404
rect 33508 13184 33560 13190
rect 33508 13126 33560 13132
rect 33416 12980 33468 12986
rect 33416 12922 33468 12928
rect 33322 12336 33378 12345
rect 33322 12271 33324 12280
rect 33376 12271 33378 12280
rect 33324 12242 33376 12248
rect 33152 11614 33272 11642
rect 32956 11348 33008 11354
rect 32956 11290 33008 11296
rect 33048 11212 33100 11218
rect 33048 11154 33100 11160
rect 32956 11076 33008 11082
rect 32956 11018 33008 11024
rect 32968 9761 32996 11018
rect 33060 10742 33088 11154
rect 33048 10736 33100 10742
rect 33048 10678 33100 10684
rect 33152 10266 33180 11614
rect 33232 11552 33284 11558
rect 33232 11494 33284 11500
rect 33140 10260 33192 10266
rect 33140 10202 33192 10208
rect 33244 10062 33272 11494
rect 33336 10985 33364 12242
rect 33416 12232 33468 12238
rect 33416 12174 33468 12180
rect 33428 11898 33456 12174
rect 33416 11892 33468 11898
rect 33416 11834 33468 11840
rect 33520 11778 33548 13126
rect 33612 12850 33640 13398
rect 33600 12844 33652 12850
rect 33600 12786 33652 12792
rect 33704 12356 33732 14010
rect 33888 13938 33916 14214
rect 33876 13932 33928 13938
rect 33876 13874 33928 13880
rect 33888 13530 33916 13874
rect 33876 13524 33928 13530
rect 33876 13466 33928 13472
rect 33980 13326 34008 14214
rect 33968 13320 34020 13326
rect 33968 13262 34020 13268
rect 34244 13320 34296 13326
rect 34244 13262 34296 13268
rect 34256 12986 34284 13262
rect 34348 13190 34376 14962
rect 34440 14278 34468 15030
rect 34428 14272 34480 14278
rect 34428 14214 34480 14220
rect 34520 13932 34572 13938
rect 34520 13874 34572 13880
rect 34336 13184 34388 13190
rect 34336 13126 34388 13132
rect 34532 12986 34560 13874
rect 34244 12980 34296 12986
rect 34244 12922 34296 12928
rect 34520 12980 34572 12986
rect 34520 12922 34572 12928
rect 33968 12844 34020 12850
rect 33968 12786 34020 12792
rect 34336 12844 34388 12850
rect 34336 12786 34388 12792
rect 33428 11750 33548 11778
rect 33612 12328 33732 12356
rect 33322 10976 33378 10985
rect 33322 10911 33378 10920
rect 33232 10056 33284 10062
rect 33232 9998 33284 10004
rect 32954 9752 33010 9761
rect 32954 9687 33010 9696
rect 33244 9674 33272 9998
rect 33322 9752 33378 9761
rect 33322 9687 33378 9696
rect 33152 9646 33272 9674
rect 32956 9614 33008 9620
rect 32956 9556 33008 9562
rect 33048 9580 33100 9586
rect 32968 9330 32996 9556
rect 33048 9522 33100 9528
rect 33060 9489 33088 9522
rect 33046 9480 33102 9489
rect 33152 9450 33180 9646
rect 33336 9586 33364 9687
rect 33324 9580 33376 9586
rect 33324 9522 33376 9528
rect 33046 9415 33102 9424
rect 33140 9444 33192 9450
rect 33140 9386 33192 9392
rect 32968 9302 33180 9330
rect 32864 9172 32916 9178
rect 32864 9114 32916 9120
rect 33048 9172 33100 9178
rect 33048 9114 33100 9120
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 32770 8800 32826 8809
rect 32770 8735 32826 8744
rect 32864 8560 32916 8566
rect 32864 8502 32916 8508
rect 32876 8430 32904 8502
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 32864 8424 32916 8430
rect 32864 8366 32916 8372
rect 32784 8129 32812 8366
rect 32770 8120 32826 8129
rect 32968 8090 32996 8910
rect 32770 8055 32826 8064
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 32772 8016 32824 8022
rect 32772 7958 32824 7964
rect 32784 7342 32812 7958
rect 32864 7472 32916 7478
rect 32864 7414 32916 7420
rect 32680 7336 32732 7342
rect 32680 7278 32732 7284
rect 32772 7336 32824 7342
rect 32772 7278 32824 7284
rect 32692 6882 32720 7278
rect 32692 6854 32812 6882
rect 32680 6792 32732 6798
rect 32680 6734 32732 6740
rect 32588 6452 32640 6458
rect 32588 6394 32640 6400
rect 32692 6390 32720 6734
rect 32680 6384 32732 6390
rect 32680 6326 32732 6332
rect 32586 6216 32642 6225
rect 32586 6151 32642 6160
rect 32600 5778 32628 6151
rect 32588 5772 32640 5778
rect 32588 5714 32640 5720
rect 32496 5296 32548 5302
rect 32496 5238 32548 5244
rect 32508 4826 32536 5238
rect 32692 5234 32720 6326
rect 32680 5228 32732 5234
rect 32680 5170 32732 5176
rect 32784 5098 32812 6854
rect 32772 5092 32824 5098
rect 32772 5034 32824 5040
rect 32496 4820 32548 4826
rect 32496 4762 32548 4768
rect 32784 4282 32812 5034
rect 32876 4622 32904 7414
rect 32968 5846 32996 8026
rect 32956 5840 33008 5846
rect 32956 5782 33008 5788
rect 33060 5642 33088 9114
rect 33152 8022 33180 9302
rect 33232 8492 33284 8498
rect 33232 8434 33284 8440
rect 33140 8016 33192 8022
rect 33140 7958 33192 7964
rect 33140 7880 33192 7886
rect 33244 7868 33272 8434
rect 33192 7840 33272 7868
rect 33140 7822 33192 7828
rect 33232 7200 33284 7206
rect 33230 7168 33232 7177
rect 33284 7168 33286 7177
rect 33230 7103 33286 7112
rect 33140 6724 33192 6730
rect 33140 6666 33192 6672
rect 33152 6390 33180 6666
rect 33140 6384 33192 6390
rect 33140 6326 33192 6332
rect 33140 6248 33192 6254
rect 33140 6190 33192 6196
rect 33152 5778 33180 6190
rect 33140 5772 33192 5778
rect 33140 5714 33192 5720
rect 33244 5642 33272 7103
rect 33048 5636 33100 5642
rect 33048 5578 33100 5584
rect 33232 5636 33284 5642
rect 33232 5578 33284 5584
rect 33060 5370 33088 5578
rect 33048 5364 33100 5370
rect 33048 5306 33100 5312
rect 33244 5166 33272 5578
rect 33428 5166 33456 11750
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 33520 11286 33548 11630
rect 33508 11280 33560 11286
rect 33508 11222 33560 11228
rect 33508 9988 33560 9994
rect 33508 9930 33560 9936
rect 33520 9450 33548 9930
rect 33508 9444 33560 9450
rect 33508 9386 33560 9392
rect 33612 9178 33640 12328
rect 33692 12232 33744 12238
rect 33692 12174 33744 12180
rect 33876 12232 33928 12238
rect 33980 12209 34008 12786
rect 34152 12640 34204 12646
rect 34152 12582 34204 12588
rect 33876 12174 33928 12180
rect 33966 12200 34022 12209
rect 33704 10810 33732 12174
rect 33784 12164 33836 12170
rect 33784 12106 33836 12112
rect 33796 11898 33824 12106
rect 33784 11892 33836 11898
rect 33784 11834 33836 11840
rect 33888 11830 33916 12174
rect 33966 12135 34022 12144
rect 34060 12164 34112 12170
rect 34060 12106 34112 12112
rect 34072 12050 34100 12106
rect 33980 12022 34100 12050
rect 33876 11824 33928 11830
rect 33876 11766 33928 11772
rect 33980 11762 34008 12022
rect 34060 11892 34112 11898
rect 34060 11834 34112 11840
rect 33968 11756 34020 11762
rect 33968 11698 34020 11704
rect 33980 11558 34008 11698
rect 33968 11552 34020 11558
rect 33968 11494 34020 11500
rect 33782 11384 33838 11393
rect 33782 11319 33784 11328
rect 33836 11319 33838 11328
rect 33968 11348 34020 11354
rect 33784 11290 33836 11296
rect 33968 11290 34020 11296
rect 33692 10804 33744 10810
rect 33692 10746 33744 10752
rect 33876 10668 33928 10674
rect 33876 10610 33928 10616
rect 33784 10260 33836 10266
rect 33784 10202 33836 10208
rect 33690 10024 33746 10033
rect 33690 9959 33692 9968
rect 33744 9959 33746 9968
rect 33692 9930 33744 9936
rect 33600 9172 33652 9178
rect 33600 9114 33652 9120
rect 33600 8968 33652 8974
rect 33600 8910 33652 8916
rect 33612 8498 33640 8910
rect 33600 8492 33652 8498
rect 33600 8434 33652 8440
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 33600 8288 33652 8294
rect 33600 8230 33652 8236
rect 33612 7886 33640 8230
rect 33704 8090 33732 8366
rect 33692 8084 33744 8090
rect 33692 8026 33744 8032
rect 33600 7880 33652 7886
rect 33600 7822 33652 7828
rect 33796 7410 33824 10202
rect 33888 10130 33916 10610
rect 33980 10130 34008 11290
rect 34072 10180 34100 11834
rect 34164 10305 34192 12582
rect 34348 11830 34376 12786
rect 34428 12300 34480 12306
rect 34428 12242 34480 12248
rect 34336 11824 34388 11830
rect 34336 11766 34388 11772
rect 34244 11756 34296 11762
rect 34244 11698 34296 11704
rect 34256 11082 34284 11698
rect 34440 11150 34468 12242
rect 34428 11144 34480 11150
rect 34428 11086 34480 11092
rect 34244 11076 34296 11082
rect 34244 11018 34296 11024
rect 34256 10606 34284 11018
rect 34244 10600 34296 10606
rect 34242 10568 34244 10577
rect 34336 10600 34388 10606
rect 34296 10568 34298 10577
rect 34336 10542 34388 10548
rect 34242 10503 34298 10512
rect 34150 10296 34206 10305
rect 34150 10231 34206 10240
rect 34072 10152 34284 10180
rect 33876 10124 33928 10130
rect 33876 10066 33928 10072
rect 33968 10124 34020 10130
rect 33968 10066 34020 10072
rect 33888 9722 33916 10066
rect 34060 10056 34112 10062
rect 34060 9998 34112 10004
rect 34072 9761 34100 9998
rect 34150 9888 34206 9897
rect 34150 9823 34206 9832
rect 34058 9752 34114 9761
rect 33876 9716 33928 9722
rect 34058 9687 34114 9696
rect 33876 9658 33928 9664
rect 34060 9648 34112 9654
rect 34060 9590 34112 9596
rect 33876 9580 33928 9586
rect 33876 9522 33928 9528
rect 33888 9178 33916 9522
rect 34072 9382 34100 9590
rect 34060 9376 34112 9382
rect 34060 9318 34112 9324
rect 33876 9172 33928 9178
rect 33876 9114 33928 9120
rect 33600 7404 33652 7410
rect 33600 7346 33652 7352
rect 33784 7404 33836 7410
rect 33784 7346 33836 7352
rect 33508 7200 33560 7206
rect 33508 7142 33560 7148
rect 33520 6798 33548 7142
rect 33612 6934 33640 7346
rect 33692 7268 33744 7274
rect 33692 7210 33744 7216
rect 33600 6928 33652 6934
rect 33600 6870 33652 6876
rect 33508 6792 33560 6798
rect 33508 6734 33560 6740
rect 33600 6792 33652 6798
rect 33600 6734 33652 6740
rect 33506 6624 33562 6633
rect 33506 6559 33562 6568
rect 33520 6390 33548 6559
rect 33508 6384 33560 6390
rect 33508 6326 33560 6332
rect 33232 5160 33284 5166
rect 33232 5102 33284 5108
rect 33416 5160 33468 5166
rect 33416 5102 33468 5108
rect 33048 4820 33100 4826
rect 33048 4762 33100 4768
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 32772 4276 32824 4282
rect 32772 4218 32824 4224
rect 32404 4208 32456 4214
rect 32404 4150 32456 4156
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 32680 4140 32732 4146
rect 32680 4082 32732 4088
rect 32508 3534 32536 4082
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 32600 3534 32628 4014
rect 32692 3670 32720 4082
rect 32680 3664 32732 3670
rect 32680 3606 32732 3612
rect 32496 3528 32548 3534
rect 32496 3470 32548 3476
rect 32588 3528 32640 3534
rect 32588 3470 32640 3476
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 31300 2644 31352 2650
rect 31300 2586 31352 2592
rect 5540 2440 5592 2446
rect 5460 2388 5540 2394
rect 5460 2382 5592 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 31208 2440 31260 2446
rect 31208 2382 31260 2388
rect 5460 2366 5580 2382
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 32 800 60 2246
rect 5184 870 5304 898
rect 5184 800 5212 870
rect 18 200 74 800
rect 5170 200 5226 800
rect 5276 762 5304 870
rect 5460 762 5488 2366
rect 31312 2310 31340 2586
rect 32508 2582 32536 3470
rect 32680 3120 32732 3126
rect 32784 3108 32812 4218
rect 32876 3670 32904 4558
rect 33060 3942 33088 4762
rect 33428 4690 33456 5102
rect 33416 4684 33468 4690
rect 33416 4626 33468 4632
rect 33048 3936 33100 3942
rect 33048 3878 33100 3884
rect 32864 3664 32916 3670
rect 32864 3606 32916 3612
rect 32876 3126 32904 3606
rect 32732 3080 32812 3108
rect 32864 3120 32916 3126
rect 32680 3062 32732 3068
rect 32864 3062 32916 3068
rect 32496 2576 32548 2582
rect 32496 2518 32548 2524
rect 32692 2446 32720 3062
rect 33060 2774 33088 3878
rect 33612 3466 33640 6734
rect 33704 6474 33732 7210
rect 33796 6633 33824 7346
rect 33888 6798 33916 9114
rect 34164 8974 34192 9823
rect 34152 8968 34204 8974
rect 34152 8910 34204 8916
rect 34152 8424 34204 8430
rect 34152 8366 34204 8372
rect 34060 7880 34112 7886
rect 34164 7857 34192 8366
rect 34060 7822 34112 7828
rect 34150 7848 34206 7857
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 33980 6746 34008 7346
rect 34072 7002 34100 7822
rect 34150 7783 34206 7792
rect 34152 7268 34204 7274
rect 34152 7210 34204 7216
rect 34164 7002 34192 7210
rect 34060 6996 34112 7002
rect 34060 6938 34112 6944
rect 34152 6996 34204 7002
rect 34152 6938 34204 6944
rect 34072 6866 34100 6938
rect 34256 6866 34284 10152
rect 34348 10130 34376 10542
rect 34336 10124 34388 10130
rect 34336 10066 34388 10072
rect 34336 9920 34388 9926
rect 34336 9862 34388 9868
rect 34348 8838 34376 9862
rect 34440 9450 34468 11086
rect 34428 9444 34480 9450
rect 34428 9386 34480 9392
rect 34336 8832 34388 8838
rect 34336 8774 34388 8780
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 34244 6860 34296 6866
rect 34244 6802 34296 6808
rect 33980 6718 34192 6746
rect 33782 6624 33838 6633
rect 33782 6559 33838 6568
rect 33704 6446 34008 6474
rect 33980 6440 34008 6446
rect 34060 6452 34112 6458
rect 33980 6412 34060 6440
rect 34060 6394 34112 6400
rect 33692 6316 33744 6322
rect 33692 6258 33744 6264
rect 33704 4826 33732 6258
rect 33968 6112 34020 6118
rect 33968 6054 34020 6060
rect 33782 5400 33838 5409
rect 33782 5335 33784 5344
rect 33836 5335 33838 5344
rect 33784 5306 33836 5312
rect 33874 4992 33930 5001
rect 33874 4927 33930 4936
rect 33692 4820 33744 4826
rect 33692 4762 33744 4768
rect 33888 4690 33916 4927
rect 33784 4684 33836 4690
rect 33784 4626 33836 4632
rect 33876 4684 33928 4690
rect 33876 4626 33928 4632
rect 33692 3732 33744 3738
rect 33692 3674 33744 3680
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 33704 2854 33732 3674
rect 33692 2848 33744 2854
rect 33692 2790 33744 2796
rect 33796 2774 33824 4626
rect 33888 4486 33916 4626
rect 33876 4480 33928 4486
rect 33876 4422 33928 4428
rect 33876 4276 33928 4282
rect 33876 4218 33928 4224
rect 33888 4010 33916 4218
rect 33980 4146 34008 6054
rect 34072 5914 34100 6394
rect 34164 6225 34192 6718
rect 34244 6316 34296 6322
rect 34244 6258 34296 6264
rect 34150 6216 34206 6225
rect 34150 6151 34206 6160
rect 34060 5908 34112 5914
rect 34060 5850 34112 5856
rect 34256 5710 34284 6258
rect 34244 5704 34296 5710
rect 34244 5646 34296 5652
rect 34348 5137 34376 8774
rect 34440 8480 34468 9386
rect 34532 8786 34560 12922
rect 34624 10810 34652 17070
rect 34716 16522 34744 17138
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34704 16516 34756 16522
rect 34704 16458 34756 16464
rect 34716 16250 34744 16458
rect 34704 16244 34756 16250
rect 34704 16186 34756 16192
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 35624 16040 35676 16046
rect 35624 15982 35676 15988
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15428 34848 15434
rect 34796 15370 34848 15376
rect 34704 15360 34756 15366
rect 34704 15302 34756 15308
rect 34716 14822 34744 15302
rect 34704 14816 34756 14822
rect 34704 14758 34756 14764
rect 34716 13938 34744 14758
rect 34704 13932 34756 13938
rect 34704 13874 34756 13880
rect 34808 11642 34836 15370
rect 35348 15020 35400 15026
rect 35348 14962 35400 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14482 35388 14962
rect 35452 14618 35480 15982
rect 35636 15706 35664 15982
rect 35624 15700 35676 15706
rect 35624 15642 35676 15648
rect 35624 14952 35676 14958
rect 35624 14894 35676 14900
rect 35440 14612 35492 14618
rect 35440 14554 35492 14560
rect 35348 14476 35400 14482
rect 35348 14418 35400 14424
rect 34888 14408 34940 14414
rect 34888 14350 34940 14356
rect 34900 14113 34928 14350
rect 34886 14104 34942 14113
rect 34886 14039 34942 14048
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35452 13326 35480 13874
rect 35440 13320 35492 13326
rect 35440 13262 35492 13268
rect 35164 13252 35216 13258
rect 35164 13194 35216 13200
rect 35176 12850 35204 13194
rect 35348 12980 35400 12986
rect 35348 12922 35400 12928
rect 34980 12844 35032 12850
rect 34980 12786 35032 12792
rect 35164 12844 35216 12850
rect 35164 12786 35216 12792
rect 34992 12753 35020 12786
rect 35360 12782 35388 12922
rect 35348 12776 35400 12782
rect 34978 12744 35034 12753
rect 35348 12718 35400 12724
rect 34978 12679 35034 12688
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35072 12232 35124 12238
rect 35072 12174 35124 12180
rect 34888 12096 34940 12102
rect 35084 12084 35112 12174
rect 34940 12056 35112 12084
rect 35256 12096 35308 12102
rect 34888 12038 34940 12044
rect 35256 12038 35308 12044
rect 35268 11830 35296 12038
rect 35256 11824 35308 11830
rect 35256 11766 35308 11772
rect 34716 11614 34836 11642
rect 34612 10804 34664 10810
rect 34612 10746 34664 10752
rect 34612 10668 34664 10674
rect 34612 10610 34664 10616
rect 34624 9926 34652 10610
rect 34612 9920 34664 9926
rect 34612 9862 34664 9868
rect 34612 9376 34664 9382
rect 34612 9318 34664 9324
rect 34624 8974 34652 9318
rect 34612 8968 34664 8974
rect 34612 8910 34664 8916
rect 34532 8758 34652 8786
rect 34520 8492 34572 8498
rect 34440 8452 34520 8480
rect 34520 8434 34572 8440
rect 34532 8129 34560 8434
rect 34624 8362 34652 8758
rect 34716 8430 34744 11614
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34888 11280 34940 11286
rect 34888 11222 34940 11228
rect 34900 10554 34928 11222
rect 35360 10810 35388 11494
rect 35452 11014 35480 13262
rect 35636 11914 35664 14894
rect 35728 14074 35756 20946
rect 35992 20392 36044 20398
rect 35992 20334 36044 20340
rect 35808 19848 35860 19854
rect 35808 19790 35860 19796
rect 35820 18834 35848 19790
rect 35808 18828 35860 18834
rect 35808 18770 35860 18776
rect 36004 18766 36032 20334
rect 36084 20256 36136 20262
rect 36082 20224 36084 20233
rect 36136 20224 36138 20233
rect 36082 20159 36138 20168
rect 36096 19786 36124 20159
rect 36084 19780 36136 19786
rect 36084 19722 36136 19728
rect 36360 19440 36412 19446
rect 36360 19382 36412 19388
rect 35992 18760 36044 18766
rect 35992 18702 36044 18708
rect 35900 15496 35952 15502
rect 35900 15438 35952 15444
rect 35808 14884 35860 14890
rect 35808 14826 35860 14832
rect 35716 14068 35768 14074
rect 35716 14010 35768 14016
rect 35820 13938 35848 14826
rect 35808 13932 35860 13938
rect 35808 13874 35860 13880
rect 35912 12986 35940 15438
rect 35900 12980 35952 12986
rect 35900 12922 35952 12928
rect 35716 12844 35768 12850
rect 35716 12786 35768 12792
rect 35900 12844 35952 12850
rect 35900 12786 35952 12792
rect 35544 11886 35664 11914
rect 35544 11150 35572 11886
rect 35624 11756 35676 11762
rect 35624 11698 35676 11704
rect 35636 11354 35664 11698
rect 35624 11348 35676 11354
rect 35624 11290 35676 11296
rect 35624 11212 35676 11218
rect 35624 11154 35676 11160
rect 35532 11144 35584 11150
rect 35636 11121 35664 11154
rect 35532 11086 35584 11092
rect 35622 11112 35678 11121
rect 35440 11008 35492 11014
rect 35440 10950 35492 10956
rect 35348 10804 35400 10810
rect 35348 10746 35400 10752
rect 34808 10526 34928 10554
rect 35256 10600 35308 10606
rect 35256 10542 35308 10548
rect 34808 9926 34836 10526
rect 35268 10418 35296 10542
rect 35268 10390 35388 10418
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34796 9920 34848 9926
rect 34796 9862 34848 9868
rect 34808 9178 34836 9862
rect 35360 9382 35388 10390
rect 35452 9518 35480 10950
rect 35544 10470 35572 11086
rect 35622 11047 35678 11056
rect 35532 10464 35584 10470
rect 35532 10406 35584 10412
rect 35440 9512 35492 9518
rect 35440 9454 35492 9460
rect 35348 9376 35400 9382
rect 35348 9318 35400 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 9172 34848 9178
rect 34796 9114 34848 9120
rect 35072 9172 35124 9178
rect 35072 9114 35124 9120
rect 35084 8974 35112 9114
rect 35256 9036 35308 9042
rect 35256 8978 35308 8984
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 35072 8968 35124 8974
rect 35072 8910 35124 8916
rect 34704 8424 34756 8430
rect 34704 8366 34756 8372
rect 34612 8356 34664 8362
rect 34612 8298 34664 8304
rect 34518 8120 34574 8129
rect 34624 8090 34652 8298
rect 34518 8055 34574 8064
rect 34612 8084 34664 8090
rect 34612 8026 34664 8032
rect 34808 7002 34836 8910
rect 34980 8832 35032 8838
rect 34980 8774 35032 8780
rect 34992 8566 35020 8774
rect 34980 8560 35032 8566
rect 35268 8537 35296 8978
rect 35348 8968 35400 8974
rect 35348 8910 35400 8916
rect 34980 8502 35032 8508
rect 35254 8528 35310 8537
rect 35254 8463 35256 8472
rect 35308 8463 35310 8472
rect 35256 8434 35308 8440
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35162 7984 35218 7993
rect 35162 7919 35164 7928
rect 35216 7919 35218 7928
rect 35164 7890 35216 7896
rect 35360 7546 35388 8910
rect 35440 8492 35492 8498
rect 35440 8434 35492 8440
rect 35452 8090 35480 8434
rect 35544 8362 35572 10406
rect 35636 8786 35664 11047
rect 35728 9178 35756 12786
rect 35912 12102 35940 12786
rect 35900 12096 35952 12102
rect 35900 12038 35952 12044
rect 35808 11892 35860 11898
rect 35808 11834 35860 11840
rect 35820 11286 35848 11834
rect 35900 11348 35952 11354
rect 35900 11290 35952 11296
rect 35808 11280 35860 11286
rect 35808 11222 35860 11228
rect 35912 10606 35940 11290
rect 35900 10600 35952 10606
rect 35900 10542 35952 10548
rect 36004 10198 36032 18702
rect 36268 17128 36320 17134
rect 36268 17070 36320 17076
rect 36280 15706 36308 17070
rect 36268 15700 36320 15706
rect 36268 15642 36320 15648
rect 36372 15570 36400 19382
rect 36464 17882 36492 23122
rect 37280 23112 37332 23118
rect 37280 23054 37332 23060
rect 36728 23044 36780 23050
rect 36728 22986 36780 22992
rect 36740 21690 36768 22986
rect 37292 22710 37320 23054
rect 37280 22704 37332 22710
rect 37280 22646 37332 22652
rect 37476 22642 37504 23122
rect 37752 22778 37780 24550
rect 38028 24206 38056 25230
rect 38212 24954 38240 25230
rect 38200 24948 38252 24954
rect 38200 24890 38252 24896
rect 38384 24812 38436 24818
rect 38384 24754 38436 24760
rect 38396 24410 38424 24754
rect 38384 24404 38436 24410
rect 38384 24346 38436 24352
rect 38488 24206 38516 26250
rect 38936 26240 38988 26246
rect 38936 26182 38988 26188
rect 38948 25906 38976 26182
rect 38936 25900 38988 25906
rect 38936 25842 38988 25848
rect 39028 25900 39080 25906
rect 39028 25842 39080 25848
rect 39040 25362 39068 25842
rect 39028 25356 39080 25362
rect 39028 25298 39080 25304
rect 40052 25294 40080 26454
rect 40420 25498 40448 56782
rect 40408 25492 40460 25498
rect 40408 25434 40460 25440
rect 38844 25288 38896 25294
rect 38844 25230 38896 25236
rect 39212 25288 39264 25294
rect 39212 25230 39264 25236
rect 39396 25288 39448 25294
rect 39396 25230 39448 25236
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 40224 25288 40276 25294
rect 40224 25230 40276 25236
rect 38856 24682 38884 25230
rect 38844 24676 38896 24682
rect 38844 24618 38896 24624
rect 38752 24268 38804 24274
rect 38752 24210 38804 24216
rect 38016 24200 38068 24206
rect 38016 24142 38068 24148
rect 38476 24200 38528 24206
rect 38476 24142 38528 24148
rect 38488 23798 38516 24142
rect 38764 23866 38792 24210
rect 39224 24070 39252 25230
rect 39408 24682 39436 25230
rect 39948 24812 40000 24818
rect 39948 24754 40000 24760
rect 39396 24676 39448 24682
rect 39396 24618 39448 24624
rect 39212 24064 39264 24070
rect 39212 24006 39264 24012
rect 39960 23866 39988 24754
rect 40052 24750 40080 25230
rect 40236 24954 40264 25230
rect 40224 24948 40276 24954
rect 40224 24890 40276 24896
rect 40316 24812 40368 24818
rect 40316 24754 40368 24760
rect 40040 24744 40092 24750
rect 40040 24686 40092 24692
rect 40052 24410 40080 24686
rect 40040 24404 40092 24410
rect 40040 24346 40092 24352
rect 40328 24274 40356 24754
rect 40316 24268 40368 24274
rect 40316 24210 40368 24216
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 40592 24200 40644 24206
rect 40592 24142 40644 24148
rect 43444 24200 43496 24206
rect 43444 24142 43496 24148
rect 38752 23860 38804 23866
rect 38752 23802 38804 23808
rect 39948 23860 40000 23866
rect 39948 23802 40000 23808
rect 38476 23792 38528 23798
rect 38476 23734 38528 23740
rect 38488 23322 38516 23734
rect 39120 23724 39172 23730
rect 39120 23666 39172 23672
rect 39132 23322 39160 23666
rect 40144 23662 40172 24142
rect 40224 24064 40276 24070
rect 40224 24006 40276 24012
rect 40236 23866 40264 24006
rect 40224 23860 40276 23866
rect 40224 23802 40276 23808
rect 40236 23730 40264 23802
rect 40604 23730 40632 24142
rect 41236 24132 41288 24138
rect 41236 24074 41288 24080
rect 41248 23730 41276 24074
rect 42892 23860 42944 23866
rect 42892 23802 42944 23808
rect 40224 23724 40276 23730
rect 40224 23666 40276 23672
rect 40592 23724 40644 23730
rect 40592 23666 40644 23672
rect 41236 23724 41288 23730
rect 41236 23666 41288 23672
rect 40132 23656 40184 23662
rect 40132 23598 40184 23604
rect 38476 23316 38528 23322
rect 38476 23258 38528 23264
rect 39120 23316 39172 23322
rect 39120 23258 39172 23264
rect 38108 23112 38160 23118
rect 38108 23054 38160 23060
rect 38292 23112 38344 23118
rect 38292 23054 38344 23060
rect 38120 22982 38148 23054
rect 38108 22976 38160 22982
rect 38108 22918 38160 22924
rect 37740 22772 37792 22778
rect 37740 22714 37792 22720
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 36728 21684 36780 21690
rect 36728 21626 36780 21632
rect 36636 21548 36688 21554
rect 36636 21490 36688 21496
rect 37372 21548 37424 21554
rect 37372 21490 37424 21496
rect 36648 20806 36676 21490
rect 37384 20942 37412 21490
rect 37556 21480 37608 21486
rect 37556 21422 37608 21428
rect 37568 20942 37596 21422
rect 38120 21146 38148 22918
rect 38200 21548 38252 21554
rect 38200 21490 38252 21496
rect 38108 21140 38160 21146
rect 38108 21082 38160 21088
rect 38212 21010 38240 21490
rect 38304 21146 38332 23054
rect 39028 22704 39080 22710
rect 39028 22646 39080 22652
rect 38936 22092 38988 22098
rect 38936 22034 38988 22040
rect 38948 21894 38976 22034
rect 39040 22030 39068 22646
rect 40144 22642 40172 23598
rect 39212 22636 39264 22642
rect 39212 22578 39264 22584
rect 40132 22636 40184 22642
rect 40132 22578 40184 22584
rect 39120 22500 39172 22506
rect 39120 22442 39172 22448
rect 39028 22024 39080 22030
rect 39028 21966 39080 21972
rect 38936 21888 38988 21894
rect 38936 21830 38988 21836
rect 38476 21480 38528 21486
rect 38476 21422 38528 21428
rect 38292 21140 38344 21146
rect 38292 21082 38344 21088
rect 38200 21004 38252 21010
rect 38200 20946 38252 20952
rect 38488 20942 38516 21422
rect 37372 20936 37424 20942
rect 37372 20878 37424 20884
rect 37556 20936 37608 20942
rect 37556 20878 37608 20884
rect 38476 20936 38528 20942
rect 38476 20878 38528 20884
rect 36636 20800 36688 20806
rect 36636 20742 36688 20748
rect 36728 20460 36780 20466
rect 36912 20460 36964 20466
rect 36780 20420 36860 20448
rect 36728 20402 36780 20408
rect 36728 20256 36780 20262
rect 36728 20198 36780 20204
rect 36740 19922 36768 20198
rect 36544 19916 36596 19922
rect 36544 19858 36596 19864
rect 36728 19916 36780 19922
rect 36728 19858 36780 19864
rect 36556 19242 36584 19858
rect 36832 19718 36860 20420
rect 36912 20402 36964 20408
rect 36820 19712 36872 19718
rect 36820 19654 36872 19660
rect 36544 19236 36596 19242
rect 36544 19178 36596 19184
rect 36728 19236 36780 19242
rect 36728 19178 36780 19184
rect 36556 18290 36584 19178
rect 36740 18766 36768 19178
rect 36728 18760 36780 18766
rect 36728 18702 36780 18708
rect 36636 18624 36688 18630
rect 36636 18566 36688 18572
rect 36728 18624 36780 18630
rect 36728 18566 36780 18572
rect 36648 18290 36676 18566
rect 36740 18426 36768 18566
rect 36728 18420 36780 18426
rect 36728 18362 36780 18368
rect 36544 18284 36596 18290
rect 36544 18226 36596 18232
rect 36636 18284 36688 18290
rect 36636 18226 36688 18232
rect 36452 17876 36504 17882
rect 36452 17818 36504 17824
rect 36648 17678 36676 18226
rect 36728 18216 36780 18222
rect 36728 18158 36780 18164
rect 36636 17672 36688 17678
rect 36636 17614 36688 17620
rect 36648 17542 36676 17614
rect 36636 17536 36688 17542
rect 36636 17478 36688 17484
rect 36648 16590 36676 17478
rect 36636 16584 36688 16590
rect 36636 16526 36688 16532
rect 36740 16114 36768 18158
rect 36832 16250 36860 19654
rect 36924 19514 36952 20402
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 36912 19508 36964 19514
rect 36912 19450 36964 19456
rect 36912 18760 36964 18766
rect 36912 18702 36964 18708
rect 36924 18086 36952 18702
rect 37372 18624 37424 18630
rect 37372 18566 37424 18572
rect 37384 18358 37412 18566
rect 37372 18352 37424 18358
rect 37372 18294 37424 18300
rect 37476 18222 37504 19790
rect 37568 18970 37596 20878
rect 38016 19916 38068 19922
rect 38016 19858 38068 19864
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37844 19378 37872 19790
rect 38028 19378 38056 19858
rect 37832 19372 37884 19378
rect 37832 19314 37884 19320
rect 38016 19372 38068 19378
rect 38016 19314 38068 19320
rect 37556 18964 37608 18970
rect 37556 18906 37608 18912
rect 37832 18692 37884 18698
rect 37832 18634 37884 18640
rect 37464 18216 37516 18222
rect 37464 18158 37516 18164
rect 36912 18080 36964 18086
rect 36912 18022 36964 18028
rect 37372 18080 37424 18086
rect 37372 18022 37424 18028
rect 37188 17672 37240 17678
rect 37188 17614 37240 17620
rect 37280 17672 37332 17678
rect 37280 17614 37332 17620
rect 36912 17060 36964 17066
rect 36912 17002 36964 17008
rect 36924 16726 36952 17002
rect 37200 16998 37228 17614
rect 37292 17338 37320 17614
rect 37280 17332 37332 17338
rect 37280 17274 37332 17280
rect 37188 16992 37240 16998
rect 37188 16934 37240 16940
rect 36912 16720 36964 16726
rect 36912 16662 36964 16668
rect 36820 16244 36872 16250
rect 36820 16186 36872 16192
rect 36728 16108 36780 16114
rect 36728 16050 36780 16056
rect 36740 15638 36768 16050
rect 36728 15632 36780 15638
rect 36728 15574 36780 15580
rect 36360 15564 36412 15570
rect 36360 15506 36412 15512
rect 36636 15496 36688 15502
rect 36636 15438 36688 15444
rect 36360 15428 36412 15434
rect 36360 15370 36412 15376
rect 36452 15428 36504 15434
rect 36452 15370 36504 15376
rect 36176 15156 36228 15162
rect 36176 15098 36228 15104
rect 36188 14278 36216 15098
rect 36372 15026 36400 15370
rect 36360 15020 36412 15026
rect 36360 14962 36412 14968
rect 36268 14544 36320 14550
rect 36268 14486 36320 14492
rect 36176 14272 36228 14278
rect 36176 14214 36228 14220
rect 36280 13938 36308 14486
rect 36372 14482 36400 14962
rect 36360 14476 36412 14482
rect 36360 14418 36412 14424
rect 36268 13932 36320 13938
rect 36268 13874 36320 13880
rect 36084 13864 36136 13870
rect 36084 13806 36136 13812
rect 36096 12850 36124 13806
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 36084 12844 36136 12850
rect 36084 12786 36136 12792
rect 36084 12708 36136 12714
rect 36188 12696 36216 13262
rect 36280 12850 36308 13874
rect 36372 13870 36400 14418
rect 36360 13864 36412 13870
rect 36360 13806 36412 13812
rect 36464 12986 36492 15370
rect 36648 15162 36676 15438
rect 36636 15156 36688 15162
rect 36636 15098 36688 15104
rect 36544 15020 36596 15026
rect 36544 14962 36596 14968
rect 36556 14618 36584 14962
rect 36740 14634 36768 15574
rect 36544 14612 36596 14618
rect 36740 14606 36860 14634
rect 36544 14554 36596 14560
rect 36832 14550 36860 14606
rect 36820 14544 36872 14550
rect 36820 14486 36872 14492
rect 37004 14340 37056 14346
rect 37004 14282 37056 14288
rect 36728 14272 36780 14278
rect 36728 14214 36780 14220
rect 36740 13530 36768 14214
rect 37016 14074 37044 14282
rect 37004 14068 37056 14074
rect 37004 14010 37056 14016
rect 36912 13932 36964 13938
rect 36912 13874 36964 13880
rect 36728 13524 36780 13530
rect 36728 13466 36780 13472
rect 36728 13252 36780 13258
rect 36728 13194 36780 13200
rect 36820 13252 36872 13258
rect 36820 13194 36872 13200
rect 36452 12980 36504 12986
rect 36452 12922 36504 12928
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 36544 12844 36596 12850
rect 36544 12786 36596 12792
rect 36636 12844 36688 12850
rect 36636 12786 36688 12792
rect 36136 12668 36216 12696
rect 36084 12650 36136 12656
rect 36096 11762 36124 12650
rect 36360 12232 36412 12238
rect 36360 12174 36412 12180
rect 36176 12096 36228 12102
rect 36176 12038 36228 12044
rect 36084 11756 36136 11762
rect 36084 11698 36136 11704
rect 36084 11552 36136 11558
rect 36084 11494 36136 11500
rect 35992 10192 36044 10198
rect 35992 10134 36044 10140
rect 35808 10056 35860 10062
rect 35808 9998 35860 10004
rect 35820 9926 35848 9998
rect 35808 9920 35860 9926
rect 35808 9862 35860 9868
rect 35806 9480 35862 9489
rect 35806 9415 35862 9424
rect 35716 9172 35768 9178
rect 35716 9114 35768 9120
rect 35820 8906 35848 9415
rect 35808 8900 35860 8906
rect 35808 8842 35860 8848
rect 35992 8832 36044 8838
rect 35898 8800 35954 8809
rect 35636 8758 35848 8786
rect 35716 8560 35768 8566
rect 35716 8502 35768 8508
rect 35624 8492 35676 8498
rect 35624 8434 35676 8440
rect 35532 8356 35584 8362
rect 35532 8298 35584 8304
rect 35636 8090 35664 8434
rect 35440 8084 35492 8090
rect 35440 8026 35492 8032
rect 35624 8084 35676 8090
rect 35624 8026 35676 8032
rect 35622 7576 35678 7585
rect 35348 7540 35400 7546
rect 35728 7562 35756 8502
rect 35820 7970 35848 8758
rect 35954 8780 35992 8786
rect 35954 8774 36044 8780
rect 35954 8758 36032 8774
rect 35898 8735 35954 8744
rect 35912 8498 35940 8735
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 35992 8084 36044 8090
rect 35992 8026 36044 8032
rect 36004 7993 36032 8026
rect 35990 7984 36046 7993
rect 35820 7942 35940 7970
rect 35912 7886 35940 7942
rect 35990 7919 36046 7928
rect 35900 7880 35952 7886
rect 35900 7822 35952 7828
rect 35400 7500 35480 7528
rect 35678 7534 35756 7562
rect 35622 7511 35624 7520
rect 35348 7482 35400 7488
rect 35348 7336 35400 7342
rect 35348 7278 35400 7284
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6996 34848 7002
rect 34796 6938 34848 6944
rect 34704 6928 34756 6934
rect 34704 6870 34756 6876
rect 34612 6384 34664 6390
rect 34612 6326 34664 6332
rect 34428 5908 34480 5914
rect 34428 5850 34480 5856
rect 34334 5128 34390 5137
rect 34334 5063 34390 5072
rect 34152 4820 34204 4826
rect 34152 4762 34204 4768
rect 34060 4480 34112 4486
rect 34060 4422 34112 4428
rect 34072 4282 34100 4422
rect 34164 4282 34192 4762
rect 34060 4276 34112 4282
rect 34060 4218 34112 4224
rect 34152 4276 34204 4282
rect 34152 4218 34204 4224
rect 33968 4140 34020 4146
rect 33968 4082 34020 4088
rect 33876 4004 33928 4010
rect 33876 3946 33928 3952
rect 33888 3534 33916 3946
rect 33980 3602 34008 4082
rect 34152 4072 34204 4078
rect 34152 4014 34204 4020
rect 34060 3664 34112 3670
rect 34060 3606 34112 3612
rect 33968 3596 34020 3602
rect 33968 3538 34020 3544
rect 34072 3534 34100 3606
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 34060 3528 34112 3534
rect 34060 3470 34112 3476
rect 33060 2746 33180 2774
rect 33796 2746 33916 2774
rect 33152 2446 33180 2746
rect 33888 2582 33916 2746
rect 33876 2576 33928 2582
rect 33876 2518 33928 2524
rect 34164 2446 34192 4014
rect 34336 3596 34388 3602
rect 34336 3538 34388 3544
rect 34244 3460 34296 3466
rect 34244 3402 34296 3408
rect 34256 2922 34284 3402
rect 34348 3194 34376 3538
rect 34336 3188 34388 3194
rect 34336 3130 34388 3136
rect 34244 2916 34296 2922
rect 34244 2858 34296 2864
rect 32680 2440 32732 2446
rect 32680 2382 32732 2388
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 34152 2440 34204 2446
rect 34152 2382 34204 2388
rect 33508 2372 33560 2378
rect 33508 2314 33560 2320
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 22836 2304 22888 2310
rect 22836 2246 22888 2252
rect 27712 2304 27764 2310
rect 27712 2246 27764 2252
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 10980 800 11008 2246
rect 16776 800 16804 2246
rect 17696 2106 17724 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 17684 2100 17736 2106
rect 17684 2042 17736 2048
rect 21928 800 21956 2246
rect 22848 2038 22876 2246
rect 22836 2032 22888 2038
rect 22836 1974 22888 1980
rect 27724 800 27752 2246
rect 33520 800 33548 2314
rect 34440 2310 34468 5850
rect 34624 5642 34652 6326
rect 34612 5636 34664 5642
rect 34612 5578 34664 5584
rect 34520 5160 34572 5166
rect 34520 5102 34572 5108
rect 34532 3194 34560 5102
rect 34624 4758 34652 5578
rect 34716 5574 34744 6870
rect 34796 6248 34848 6254
rect 34796 6190 34848 6196
rect 34704 5568 34756 5574
rect 34704 5510 34756 5516
rect 34808 5386 34836 6190
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35360 5778 35388 7278
rect 35452 7002 35480 7500
rect 35676 7511 35678 7520
rect 35624 7482 35676 7488
rect 35716 7472 35768 7478
rect 35716 7414 35768 7420
rect 35530 7304 35586 7313
rect 35530 7239 35532 7248
rect 35584 7239 35586 7248
rect 35532 7210 35584 7216
rect 35440 6996 35492 7002
rect 35440 6938 35492 6944
rect 35624 6928 35676 6934
rect 35624 6870 35676 6876
rect 35440 6180 35492 6186
rect 35440 6122 35492 6128
rect 35164 5772 35216 5778
rect 35348 5772 35400 5778
rect 35216 5732 35296 5760
rect 35164 5714 35216 5720
rect 35268 5574 35296 5732
rect 35348 5714 35400 5720
rect 35072 5568 35124 5574
rect 35072 5510 35124 5516
rect 35256 5568 35308 5574
rect 35256 5510 35308 5516
rect 35084 5409 35112 5510
rect 34716 5358 34836 5386
rect 35070 5400 35126 5409
rect 34612 4752 34664 4758
rect 34612 4694 34664 4700
rect 34624 3398 34652 4694
rect 34716 4214 34744 5358
rect 35070 5335 35126 5344
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35348 4548 35400 4554
rect 35348 4490 35400 4496
rect 34796 4276 34848 4282
rect 34796 4218 34848 4224
rect 34704 4208 34756 4214
rect 34704 4150 34756 4156
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34520 3188 34572 3194
rect 34520 3130 34572 3136
rect 34808 3126 34836 4218
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 34808 2582 34836 3062
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2576 34848 2582
rect 34796 2518 34848 2524
rect 35360 2446 35388 4490
rect 35452 3126 35480 6122
rect 35636 5914 35664 6870
rect 35728 6866 35756 7414
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 35716 6860 35768 6866
rect 35716 6802 35768 6808
rect 35728 6322 35756 6802
rect 35912 6798 35940 7346
rect 36096 6905 36124 11494
rect 36188 9994 36216 12038
rect 36372 11354 36400 12174
rect 36556 11370 36584 12786
rect 36648 12442 36676 12786
rect 36636 12436 36688 12442
rect 36636 12378 36688 12384
rect 36740 12238 36768 13194
rect 36728 12232 36780 12238
rect 36728 12174 36780 12180
rect 36832 12102 36860 13194
rect 36636 12096 36688 12102
rect 36636 12038 36688 12044
rect 36820 12096 36872 12102
rect 36820 12038 36872 12044
rect 36648 11762 36676 12038
rect 36726 11792 36782 11801
rect 36636 11756 36688 11762
rect 36726 11727 36728 11736
rect 36636 11698 36688 11704
rect 36780 11727 36782 11736
rect 36728 11698 36780 11704
rect 36728 11552 36780 11558
rect 36728 11494 36780 11500
rect 36360 11348 36412 11354
rect 36556 11342 36676 11370
rect 36360 11290 36412 11296
rect 36544 11280 36596 11286
rect 36544 11222 36596 11228
rect 36360 10736 36412 10742
rect 36360 10678 36412 10684
rect 36176 9988 36228 9994
rect 36176 9930 36228 9936
rect 36188 9654 36216 9930
rect 36176 9648 36228 9654
rect 36176 9590 36228 9596
rect 36176 9376 36228 9382
rect 36372 9364 36400 10678
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36464 10266 36492 10610
rect 36452 10260 36504 10266
rect 36452 10202 36504 10208
rect 36228 9336 36400 9364
rect 36176 9318 36228 9324
rect 36188 8945 36216 9318
rect 36464 9178 36492 10202
rect 36556 10130 36584 11222
rect 36544 10124 36596 10130
rect 36544 10066 36596 10072
rect 36544 9988 36596 9994
rect 36544 9930 36596 9936
rect 36556 9586 36584 9930
rect 36544 9580 36596 9586
rect 36544 9522 36596 9528
rect 36452 9172 36504 9178
rect 36452 9114 36504 9120
rect 36174 8936 36230 8945
rect 36230 8894 36308 8922
rect 36174 8871 36230 8880
rect 36176 8288 36228 8294
rect 36176 8230 36228 8236
rect 36188 7886 36216 8230
rect 36280 8090 36308 8894
rect 36268 8084 36320 8090
rect 36268 8026 36320 8032
rect 36176 7880 36228 7886
rect 36176 7822 36228 7828
rect 36556 7818 36584 9522
rect 36648 9042 36676 11342
rect 36740 10470 36768 11494
rect 36820 11144 36872 11150
rect 36924 11121 36952 13874
rect 37200 13870 37228 16934
rect 37384 16590 37412 18022
rect 37476 17678 37504 18158
rect 37740 17740 37792 17746
rect 37740 17682 37792 17688
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37752 17202 37780 17682
rect 37740 17196 37792 17202
rect 37740 17138 37792 17144
rect 37464 17128 37516 17134
rect 37464 17070 37516 17076
rect 37372 16584 37424 16590
rect 37372 16526 37424 16532
rect 37280 16448 37332 16454
rect 37280 16390 37332 16396
rect 37292 14074 37320 16390
rect 37384 15162 37412 16526
rect 37476 16522 37504 17070
rect 37464 16516 37516 16522
rect 37464 16458 37516 16464
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 37660 15706 37688 16050
rect 37648 15700 37700 15706
rect 37648 15642 37700 15648
rect 37372 15156 37424 15162
rect 37372 15098 37424 15104
rect 37752 14958 37780 17138
rect 37844 16454 37872 18634
rect 38028 18426 38056 19314
rect 38016 18420 38068 18426
rect 38016 18362 38068 18368
rect 38384 18284 38436 18290
rect 38384 18226 38436 18232
rect 38396 17066 38424 18226
rect 38384 17060 38436 17066
rect 38384 17002 38436 17008
rect 38384 16652 38436 16658
rect 38384 16594 38436 16600
rect 38016 16584 38068 16590
rect 38016 16526 38068 16532
rect 37832 16448 37884 16454
rect 37832 16390 37884 16396
rect 38028 16114 38056 16526
rect 38108 16448 38160 16454
rect 38108 16390 38160 16396
rect 38120 16250 38148 16390
rect 38108 16244 38160 16250
rect 38108 16186 38160 16192
rect 38016 16108 38068 16114
rect 38016 16050 38068 16056
rect 37832 15904 37884 15910
rect 37832 15846 37884 15852
rect 37844 15502 37872 15846
rect 37832 15496 37884 15502
rect 37832 15438 37884 15444
rect 37924 15020 37976 15026
rect 37924 14962 37976 14968
rect 37740 14952 37792 14958
rect 37740 14894 37792 14900
rect 37464 14816 37516 14822
rect 37464 14758 37516 14764
rect 37280 14068 37332 14074
rect 37280 14010 37332 14016
rect 37188 13864 37240 13870
rect 37188 13806 37240 13812
rect 37188 13524 37240 13530
rect 37188 13466 37240 13472
rect 37200 13394 37228 13466
rect 37188 13388 37240 13394
rect 37188 13330 37240 13336
rect 37200 12850 37228 13330
rect 37188 12844 37240 12850
rect 37188 12786 37240 12792
rect 37004 12776 37056 12782
rect 37002 12744 37004 12753
rect 37056 12744 37058 12753
rect 37002 12679 37058 12688
rect 37188 12640 37240 12646
rect 37188 12582 37240 12588
rect 37200 12442 37228 12582
rect 37188 12436 37240 12442
rect 37188 12378 37240 12384
rect 37292 12170 37320 14010
rect 37372 14000 37424 14006
rect 37372 13942 37424 13948
rect 37384 13530 37412 13942
rect 37372 13524 37424 13530
rect 37372 13466 37424 13472
rect 37280 12164 37332 12170
rect 37280 12106 37332 12112
rect 37188 11756 37240 11762
rect 37188 11698 37240 11704
rect 37004 11688 37056 11694
rect 37004 11630 37056 11636
rect 36820 11086 36872 11092
rect 36910 11112 36966 11121
rect 36728 10464 36780 10470
rect 36728 10406 36780 10412
rect 36832 9353 36860 11086
rect 36910 11047 36912 11056
rect 36964 11047 36966 11056
rect 36912 11018 36964 11024
rect 36924 10987 36952 11018
rect 36912 10056 36964 10062
rect 36912 9998 36964 10004
rect 36924 9722 36952 9998
rect 37016 9994 37044 11630
rect 37200 11150 37228 11698
rect 37280 11280 37332 11286
rect 37280 11222 37332 11228
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 37004 9988 37056 9994
rect 37004 9930 37056 9936
rect 36912 9716 36964 9722
rect 36912 9658 36964 9664
rect 37004 9512 37056 9518
rect 37004 9454 37056 9460
rect 36912 9376 36964 9382
rect 36818 9344 36874 9353
rect 36912 9318 36964 9324
rect 36818 9279 36874 9288
rect 36728 9104 36780 9110
rect 36728 9046 36780 9052
rect 36636 9036 36688 9042
rect 36636 8978 36688 8984
rect 36544 7812 36596 7818
rect 36544 7754 36596 7760
rect 36556 7392 36584 7754
rect 36648 7546 36676 8978
rect 36740 8498 36768 9046
rect 36924 8974 36952 9318
rect 36912 8968 36964 8974
rect 36912 8910 36964 8916
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36728 7880 36780 7886
rect 36728 7822 36780 7828
rect 36636 7540 36688 7546
rect 36636 7482 36688 7488
rect 36636 7404 36688 7410
rect 36556 7364 36636 7392
rect 36636 7346 36688 7352
rect 36082 6896 36138 6905
rect 36082 6831 36138 6840
rect 36450 6896 36506 6905
rect 36450 6831 36506 6840
rect 35900 6792 35952 6798
rect 35900 6734 35952 6740
rect 36084 6792 36136 6798
rect 36084 6734 36136 6740
rect 36176 6792 36228 6798
rect 36176 6734 36228 6740
rect 35716 6316 35768 6322
rect 35716 6258 35768 6264
rect 36096 6254 36124 6734
rect 36084 6248 36136 6254
rect 36084 6190 36136 6196
rect 36188 6118 36216 6734
rect 36464 6390 36492 6831
rect 36452 6384 36504 6390
rect 36452 6326 36504 6332
rect 36360 6316 36412 6322
rect 36360 6258 36412 6264
rect 36176 6112 36228 6118
rect 36176 6054 36228 6060
rect 35624 5908 35676 5914
rect 35624 5850 35676 5856
rect 36188 5710 36216 6054
rect 36372 5778 36400 6258
rect 36648 6118 36676 7346
rect 36740 6730 36768 7822
rect 37016 7342 37044 9454
rect 37096 8968 37148 8974
rect 37096 8910 37148 8916
rect 37108 8634 37136 8910
rect 37096 8628 37148 8634
rect 37096 8570 37148 8576
rect 37004 7336 37056 7342
rect 37004 7278 37056 7284
rect 37096 7268 37148 7274
rect 37096 7210 37148 7216
rect 36728 6724 36780 6730
rect 36728 6666 36780 6672
rect 37108 6322 37136 7210
rect 37200 6866 37228 11086
rect 37292 10674 37320 11222
rect 37372 11008 37424 11014
rect 37372 10950 37424 10956
rect 37280 10668 37332 10674
rect 37280 10610 37332 10616
rect 37292 9586 37320 10610
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 37292 9489 37320 9522
rect 37278 9480 37334 9489
rect 37278 9415 37334 9424
rect 37384 8820 37412 10950
rect 37476 9178 37504 14758
rect 37936 14618 37964 14962
rect 38292 14952 38344 14958
rect 38292 14894 38344 14900
rect 38200 14816 38252 14822
rect 38200 14758 38252 14764
rect 37924 14612 37976 14618
rect 37924 14554 37976 14560
rect 37556 14408 37608 14414
rect 37556 14350 37608 14356
rect 37568 11898 37596 14350
rect 38212 14278 38240 14758
rect 38304 14396 38332 14894
rect 38396 14618 38424 16594
rect 38488 15706 38516 20878
rect 38844 20460 38896 20466
rect 38844 20402 38896 20408
rect 38752 20392 38804 20398
rect 38752 20334 38804 20340
rect 38764 19990 38792 20334
rect 38856 20058 38884 20402
rect 39040 20058 39068 21966
rect 39132 21894 39160 22442
rect 39224 22094 39252 22578
rect 39224 22066 39344 22094
rect 39316 22030 39344 22066
rect 39304 22024 39356 22030
rect 39304 21966 39356 21972
rect 39120 21888 39172 21894
rect 39120 21830 39172 21836
rect 38844 20052 38896 20058
rect 38844 19994 38896 20000
rect 39028 20052 39080 20058
rect 39028 19994 39080 20000
rect 38752 19984 38804 19990
rect 38752 19926 38804 19932
rect 39132 19514 39160 21830
rect 39316 21690 39344 21966
rect 40236 21894 40264 23666
rect 40500 23112 40552 23118
rect 40500 23054 40552 23060
rect 40512 22778 40540 23054
rect 40500 22772 40552 22778
rect 40500 22714 40552 22720
rect 40500 22636 40552 22642
rect 40500 22578 40552 22584
rect 40512 22098 40540 22578
rect 40604 22574 40632 23666
rect 40868 23520 40920 23526
rect 40868 23462 40920 23468
rect 40880 23118 40908 23462
rect 40868 23112 40920 23118
rect 40868 23054 40920 23060
rect 40776 22636 40828 22642
rect 40776 22578 40828 22584
rect 40592 22568 40644 22574
rect 40592 22510 40644 22516
rect 40788 22098 40816 22578
rect 40500 22092 40552 22098
rect 40500 22034 40552 22040
rect 40776 22092 40828 22098
rect 40776 22034 40828 22040
rect 40960 22092 41012 22098
rect 40960 22034 41012 22040
rect 40788 21962 40816 22034
rect 40776 21956 40828 21962
rect 40776 21898 40828 21904
rect 40868 21956 40920 21962
rect 40868 21898 40920 21904
rect 40224 21888 40276 21894
rect 40224 21830 40276 21836
rect 40684 21888 40736 21894
rect 40684 21830 40736 21836
rect 39304 21684 39356 21690
rect 39304 21626 39356 21632
rect 40696 21622 40724 21830
rect 40880 21690 40908 21898
rect 40868 21684 40920 21690
rect 40868 21626 40920 21632
rect 40684 21616 40736 21622
rect 40684 21558 40736 21564
rect 40592 21548 40644 21554
rect 40592 21490 40644 21496
rect 39396 20800 39448 20806
rect 39396 20742 39448 20748
rect 39120 19508 39172 19514
rect 39120 19450 39172 19456
rect 39408 19446 39436 20742
rect 40040 20460 40092 20466
rect 40040 20402 40092 20408
rect 40052 19922 40080 20402
rect 40316 20392 40368 20398
rect 40316 20334 40368 20340
rect 40040 19916 40092 19922
rect 40040 19858 40092 19864
rect 40328 19854 40356 20334
rect 40604 20058 40632 21490
rect 40592 20052 40644 20058
rect 40592 19994 40644 20000
rect 40316 19848 40368 19854
rect 40316 19790 40368 19796
rect 39396 19440 39448 19446
rect 39396 19382 39448 19388
rect 39856 19440 39908 19446
rect 39856 19382 39908 19388
rect 40040 19440 40092 19446
rect 40040 19382 40092 19388
rect 39028 18896 39080 18902
rect 39028 18838 39080 18844
rect 38660 18828 38712 18834
rect 38660 18770 38712 18776
rect 38568 17604 38620 17610
rect 38568 17546 38620 17552
rect 38580 17338 38608 17546
rect 38568 17332 38620 17338
rect 38568 17274 38620 17280
rect 38580 16590 38608 17274
rect 38568 16584 38620 16590
rect 38568 16526 38620 16532
rect 38476 15700 38528 15706
rect 38476 15642 38528 15648
rect 38672 15434 38700 18770
rect 39040 18290 39068 18838
rect 39396 18828 39448 18834
rect 39396 18770 39448 18776
rect 39212 18760 39264 18766
rect 39212 18702 39264 18708
rect 39304 18760 39356 18766
rect 39304 18702 39356 18708
rect 39028 18284 39080 18290
rect 39028 18226 39080 18232
rect 38752 17876 38804 17882
rect 38752 17818 38804 17824
rect 38764 17202 38792 17818
rect 38936 17536 38988 17542
rect 38936 17478 38988 17484
rect 38948 17202 38976 17478
rect 38752 17196 38804 17202
rect 38752 17138 38804 17144
rect 38936 17196 38988 17202
rect 38936 17138 38988 17144
rect 38764 16590 38792 17138
rect 38948 17105 38976 17138
rect 38934 17096 38990 17105
rect 39040 17066 39068 18226
rect 39224 18222 39252 18702
rect 39212 18216 39264 18222
rect 39212 18158 39264 18164
rect 39224 17882 39252 18158
rect 39316 18086 39344 18702
rect 39304 18080 39356 18086
rect 39304 18022 39356 18028
rect 39212 17876 39264 17882
rect 39212 17818 39264 17824
rect 38934 17031 38990 17040
rect 39028 17060 39080 17066
rect 39028 17002 39080 17008
rect 38752 16584 38804 16590
rect 38752 16526 38804 16532
rect 38764 16114 38792 16526
rect 38752 16108 38804 16114
rect 38752 16050 38804 16056
rect 39028 15564 39080 15570
rect 39028 15506 39080 15512
rect 38660 15428 38712 15434
rect 38660 15370 38712 15376
rect 38752 15360 38804 15366
rect 38804 15320 38884 15348
rect 38752 15302 38804 15308
rect 38856 14890 38884 15320
rect 39040 15162 39068 15506
rect 39120 15496 39172 15502
rect 39120 15438 39172 15444
rect 39028 15156 39080 15162
rect 39028 15098 39080 15104
rect 39132 15094 39160 15438
rect 39408 15366 39436 18770
rect 39580 18692 39632 18698
rect 39580 18634 39632 18640
rect 39592 18290 39620 18634
rect 39580 18284 39632 18290
rect 39580 18226 39632 18232
rect 39488 16584 39540 16590
rect 39592 16572 39620 18226
rect 39868 17542 39896 19382
rect 40052 19258 40080 19382
rect 40052 19230 40172 19258
rect 40040 19168 40092 19174
rect 40040 19110 40092 19116
rect 40052 18970 40080 19110
rect 40040 18964 40092 18970
rect 40040 18906 40092 18912
rect 40144 18834 40172 19230
rect 40224 19168 40276 19174
rect 40224 19110 40276 19116
rect 40236 18834 40264 19110
rect 40328 18970 40356 19790
rect 40972 19360 41000 22034
rect 41144 22024 41196 22030
rect 41144 21966 41196 21972
rect 41052 21480 41104 21486
rect 41156 21468 41184 21966
rect 41248 21690 41276 23666
rect 41696 23520 41748 23526
rect 41696 23462 41748 23468
rect 41972 23520 42024 23526
rect 41972 23462 42024 23468
rect 41604 23112 41656 23118
rect 41604 23054 41656 23060
rect 41328 22636 41380 22642
rect 41328 22578 41380 22584
rect 41340 21962 41368 22578
rect 41616 22574 41644 23054
rect 41708 22778 41736 23462
rect 41984 23186 42012 23462
rect 41972 23180 42024 23186
rect 41972 23122 42024 23128
rect 42432 23044 42484 23050
rect 42432 22986 42484 22992
rect 42444 22778 42472 22986
rect 41696 22772 41748 22778
rect 41696 22714 41748 22720
rect 42432 22772 42484 22778
rect 42432 22714 42484 22720
rect 41604 22568 41656 22574
rect 41604 22510 41656 22516
rect 41512 22432 41564 22438
rect 41512 22374 41564 22380
rect 41328 21956 41380 21962
rect 41328 21898 41380 21904
rect 41236 21684 41288 21690
rect 41236 21626 41288 21632
rect 41104 21440 41184 21468
rect 41052 21422 41104 21428
rect 41064 20602 41092 21422
rect 41052 20596 41104 20602
rect 41052 20538 41104 20544
rect 41236 20460 41288 20466
rect 41236 20402 41288 20408
rect 41248 19514 41276 20402
rect 41420 20256 41472 20262
rect 41420 20198 41472 20204
rect 41432 19922 41460 20198
rect 41420 19916 41472 19922
rect 41420 19858 41472 19864
rect 41524 19854 41552 22374
rect 42444 22234 42472 22714
rect 42904 22710 42932 23802
rect 43456 23798 43484 24142
rect 43444 23792 43496 23798
rect 43444 23734 43496 23740
rect 43456 23322 43484 23734
rect 43444 23316 43496 23322
rect 43444 23258 43496 23264
rect 42892 22704 42944 22710
rect 42892 22646 42944 22652
rect 42432 22228 42484 22234
rect 42432 22170 42484 22176
rect 41696 22024 41748 22030
rect 41696 21966 41748 21972
rect 41708 20466 41736 21966
rect 42156 21888 42208 21894
rect 42156 21830 42208 21836
rect 42168 21622 42196 21830
rect 42064 21616 42116 21622
rect 42064 21558 42116 21564
rect 42156 21616 42208 21622
rect 42156 21558 42208 21564
rect 41696 20460 41748 20466
rect 41696 20402 41748 20408
rect 41880 20460 41932 20466
rect 41880 20402 41932 20408
rect 41512 19848 41564 19854
rect 41512 19790 41564 19796
rect 41892 19514 41920 20402
rect 41236 19508 41288 19514
rect 41236 19450 41288 19456
rect 41880 19508 41932 19514
rect 41880 19450 41932 19456
rect 41144 19372 41196 19378
rect 40972 19332 41144 19360
rect 41144 19314 41196 19320
rect 41420 19372 41472 19378
rect 41880 19372 41932 19378
rect 41420 19314 41472 19320
rect 41800 19332 41880 19360
rect 40316 18964 40368 18970
rect 40316 18906 40368 18912
rect 40132 18828 40184 18834
rect 40132 18770 40184 18776
rect 40224 18828 40276 18834
rect 40224 18770 40276 18776
rect 40144 18426 40172 18770
rect 40592 18760 40644 18766
rect 40592 18702 40644 18708
rect 40132 18420 40184 18426
rect 40132 18362 40184 18368
rect 39856 17536 39908 17542
rect 39856 17478 39908 17484
rect 39948 17196 40000 17202
rect 39948 17138 40000 17144
rect 40040 17196 40092 17202
rect 40040 17138 40092 17144
rect 40224 17196 40276 17202
rect 40224 17138 40276 17144
rect 39540 16544 39620 16572
rect 39488 16526 39540 16532
rect 39960 16046 39988 17138
rect 40052 16454 40080 17138
rect 40236 16794 40264 17138
rect 40224 16788 40276 16794
rect 40224 16730 40276 16736
rect 40040 16448 40092 16454
rect 40040 16390 40092 16396
rect 40052 16114 40080 16390
rect 40236 16250 40264 16730
rect 40316 16584 40368 16590
rect 40316 16526 40368 16532
rect 40224 16244 40276 16250
rect 40224 16186 40276 16192
rect 40040 16108 40092 16114
rect 40040 16050 40092 16056
rect 39948 16040 40000 16046
rect 39948 15982 40000 15988
rect 39948 15428 40000 15434
rect 39948 15370 40000 15376
rect 39396 15360 39448 15366
rect 39396 15302 39448 15308
rect 39960 15094 39988 15370
rect 39120 15088 39172 15094
rect 39120 15030 39172 15036
rect 39948 15088 40000 15094
rect 39948 15030 40000 15036
rect 39132 14958 39160 15030
rect 39304 15020 39356 15026
rect 39304 14962 39356 14968
rect 39120 14952 39172 14958
rect 39120 14894 39172 14900
rect 38844 14884 38896 14890
rect 38844 14826 38896 14832
rect 38384 14612 38436 14618
rect 38384 14554 38436 14560
rect 38384 14408 38436 14414
rect 38304 14368 38384 14396
rect 38384 14350 38436 14356
rect 38660 14408 38712 14414
rect 38660 14350 38712 14356
rect 38200 14272 38252 14278
rect 38200 14214 38252 14220
rect 37924 13728 37976 13734
rect 37924 13670 37976 13676
rect 37936 12986 37964 13670
rect 38108 13524 38160 13530
rect 38108 13466 38160 13472
rect 38016 13184 38068 13190
rect 38120 13138 38148 13466
rect 38068 13132 38148 13138
rect 38016 13126 38148 13132
rect 38292 13184 38344 13190
rect 38292 13126 38344 13132
rect 38028 13110 38148 13126
rect 37924 12980 37976 12986
rect 37924 12922 37976 12928
rect 37936 12374 37964 12922
rect 38120 12434 38148 13110
rect 38304 12850 38332 13126
rect 38292 12844 38344 12850
rect 38292 12786 38344 12792
rect 38028 12406 38148 12434
rect 37924 12368 37976 12374
rect 37924 12310 37976 12316
rect 37740 12300 37792 12306
rect 37792 12260 37872 12288
rect 37740 12242 37792 12248
rect 37648 12232 37700 12238
rect 37646 12200 37648 12209
rect 37700 12200 37702 12209
rect 37646 12135 37702 12144
rect 37648 12096 37700 12102
rect 37648 12038 37700 12044
rect 37556 11892 37608 11898
rect 37556 11834 37608 11840
rect 37554 11656 37610 11665
rect 37554 11591 37556 11600
rect 37608 11591 37610 11600
rect 37556 11562 37608 11568
rect 37568 11150 37596 11562
rect 37556 11144 37608 11150
rect 37556 11086 37608 11092
rect 37660 10742 37688 12038
rect 37740 11688 37792 11694
rect 37740 11630 37792 11636
rect 37752 11354 37780 11630
rect 37740 11348 37792 11354
rect 37740 11290 37792 11296
rect 37844 10742 37872 12260
rect 37924 12232 37976 12238
rect 37924 12174 37976 12180
rect 37936 11762 37964 12174
rect 37924 11756 37976 11762
rect 37924 11698 37976 11704
rect 37924 11552 37976 11558
rect 37924 11494 37976 11500
rect 37936 11354 37964 11494
rect 37924 11348 37976 11354
rect 37924 11290 37976 11296
rect 37648 10736 37700 10742
rect 37648 10678 37700 10684
rect 37832 10736 37884 10742
rect 37832 10678 37884 10684
rect 37556 10260 37608 10266
rect 37556 10202 37608 10208
rect 37464 9172 37516 9178
rect 37464 9114 37516 9120
rect 37464 8832 37516 8838
rect 37384 8792 37464 8820
rect 37464 8774 37516 8780
rect 37280 8424 37332 8430
rect 37278 8392 37280 8401
rect 37332 8392 37334 8401
rect 37278 8327 37334 8336
rect 37372 8288 37424 8294
rect 37372 8230 37424 8236
rect 37384 7018 37412 8230
rect 37476 7478 37504 8774
rect 37568 8634 37596 10202
rect 37648 9376 37700 9382
rect 37646 9344 37648 9353
rect 37700 9344 37702 9353
rect 37646 9279 37702 9288
rect 37556 8628 37608 8634
rect 37556 8570 37608 8576
rect 37740 8492 37792 8498
rect 37740 8434 37792 8440
rect 37752 8090 37780 8434
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37648 7880 37700 7886
rect 37648 7822 37700 7828
rect 37464 7472 37516 7478
rect 37464 7414 37516 7420
rect 37476 7206 37504 7414
rect 37464 7200 37516 7206
rect 37464 7142 37516 7148
rect 37384 6990 37504 7018
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 36912 6316 36964 6322
rect 36912 6258 36964 6264
rect 37096 6316 37148 6322
rect 37096 6258 37148 6264
rect 36636 6112 36688 6118
rect 36636 6054 36688 6060
rect 36924 5846 36952 6258
rect 36912 5840 36964 5846
rect 36912 5782 36964 5788
rect 36360 5772 36412 5778
rect 37004 5772 37056 5778
rect 36412 5732 36492 5760
rect 36360 5714 36412 5720
rect 36176 5704 36228 5710
rect 36176 5646 36228 5652
rect 35716 5568 35768 5574
rect 35716 5510 35768 5516
rect 35728 5137 35756 5510
rect 35808 5296 35860 5302
rect 35808 5238 35860 5244
rect 35714 5128 35770 5137
rect 35714 5063 35770 5072
rect 35820 4282 35848 5238
rect 36082 4584 36138 4593
rect 36082 4519 36084 4528
rect 36136 4519 36138 4528
rect 36084 4490 36136 4496
rect 35808 4276 35860 4282
rect 35808 4218 35860 4224
rect 35716 3460 35768 3466
rect 35716 3402 35768 3408
rect 35728 3126 35756 3402
rect 35440 3120 35492 3126
rect 35440 3062 35492 3068
rect 35716 3120 35768 3126
rect 35716 3062 35768 3068
rect 36096 2774 36124 4490
rect 36268 3664 36320 3670
rect 36268 3606 36320 3612
rect 36280 3058 36308 3606
rect 36360 3392 36412 3398
rect 36360 3334 36412 3340
rect 36268 3052 36320 3058
rect 36268 2994 36320 3000
rect 36372 2854 36400 3334
rect 36464 2922 36492 5732
rect 37056 5732 37228 5760
rect 37004 5714 37056 5720
rect 37016 5642 37044 5714
rect 37200 5658 37228 5732
rect 37004 5636 37056 5642
rect 37200 5630 37320 5658
rect 37004 5578 37056 5584
rect 37292 5545 37320 5630
rect 37278 5536 37334 5545
rect 37278 5471 37334 5480
rect 37476 5250 37504 6990
rect 37660 6798 37688 7822
rect 37648 6792 37700 6798
rect 37648 6734 37700 6740
rect 37660 5302 37688 6734
rect 37740 6724 37792 6730
rect 37740 6666 37792 6672
rect 37108 5222 37504 5250
rect 37648 5296 37700 5302
rect 37648 5238 37700 5244
rect 37108 4690 37136 5222
rect 37188 5160 37240 5166
rect 37188 5102 37240 5108
rect 37096 4684 37148 4690
rect 37096 4626 37148 4632
rect 37096 4548 37148 4554
rect 37096 4490 37148 4496
rect 37108 4282 37136 4490
rect 37096 4276 37148 4282
rect 37096 4218 37148 4224
rect 37108 3466 37136 4218
rect 37200 3738 37228 5102
rect 37280 5024 37332 5030
rect 37280 4966 37332 4972
rect 37292 4214 37320 4966
rect 37556 4820 37608 4826
rect 37556 4762 37608 4768
rect 37464 4684 37516 4690
rect 37464 4626 37516 4632
rect 37280 4208 37332 4214
rect 37280 4150 37332 4156
rect 37476 4078 37504 4626
rect 37568 4570 37596 4762
rect 37660 4570 37688 5238
rect 37568 4542 37688 4570
rect 37280 4072 37332 4078
rect 37280 4014 37332 4020
rect 37464 4072 37516 4078
rect 37464 4014 37516 4020
rect 37188 3732 37240 3738
rect 37188 3674 37240 3680
rect 37292 3602 37320 4014
rect 37372 3936 37424 3942
rect 37372 3878 37424 3884
rect 37280 3596 37332 3602
rect 37280 3538 37332 3544
rect 37096 3460 37148 3466
rect 37096 3402 37148 3408
rect 37292 3194 37320 3538
rect 37384 3448 37412 3878
rect 37464 3460 37516 3466
rect 37384 3420 37464 3448
rect 37464 3402 37516 3408
rect 37280 3188 37332 3194
rect 37280 3130 37332 3136
rect 37292 3058 37320 3130
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 36452 2916 36504 2922
rect 36452 2858 36504 2864
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 37292 2774 37320 2994
rect 37568 2990 37596 4542
rect 37648 4480 37700 4486
rect 37648 4422 37700 4428
rect 37660 3194 37688 4422
rect 37752 4078 37780 6666
rect 37844 6100 37872 10678
rect 38028 7970 38056 12406
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 38120 12102 38148 12174
rect 38108 12096 38160 12102
rect 38108 12038 38160 12044
rect 38120 11286 38148 12038
rect 38108 11280 38160 11286
rect 38108 11222 38160 11228
rect 38396 10810 38424 14350
rect 38476 14340 38528 14346
rect 38476 14282 38528 14288
rect 38488 14006 38516 14282
rect 38672 14074 38700 14350
rect 38856 14074 38884 14826
rect 38660 14068 38712 14074
rect 38660 14010 38712 14016
rect 38844 14068 38896 14074
rect 38844 14010 38896 14016
rect 38476 14000 38528 14006
rect 38476 13942 38528 13948
rect 38488 13802 38516 13942
rect 38476 13796 38528 13802
rect 38476 13738 38528 13744
rect 38488 11694 38516 13738
rect 38660 13388 38712 13394
rect 38660 13330 38712 13336
rect 38568 13184 38620 13190
rect 38568 13126 38620 13132
rect 38580 12102 38608 13126
rect 38568 12096 38620 12102
rect 38568 12038 38620 12044
rect 38672 11762 38700 13330
rect 38856 12442 38884 14010
rect 39132 13870 39160 14894
rect 39212 14816 39264 14822
rect 39212 14758 39264 14764
rect 39224 13938 39252 14758
rect 39316 14482 39344 14962
rect 39488 14952 39540 14958
rect 39488 14894 39540 14900
rect 39500 14550 39528 14894
rect 39488 14544 39540 14550
rect 39488 14486 39540 14492
rect 39304 14476 39356 14482
rect 39304 14418 39356 14424
rect 39212 13932 39264 13938
rect 39212 13874 39264 13880
rect 39120 13864 39172 13870
rect 39120 13806 39172 13812
rect 39212 13728 39264 13734
rect 39212 13670 39264 13676
rect 39224 13530 39252 13670
rect 39212 13524 39264 13530
rect 39212 13466 39264 13472
rect 39120 13456 39172 13462
rect 39120 13398 39172 13404
rect 38936 12776 38988 12782
rect 38936 12718 38988 12724
rect 38844 12436 38896 12442
rect 38844 12378 38896 12384
rect 38660 11756 38712 11762
rect 38660 11698 38712 11704
rect 38476 11688 38528 11694
rect 38476 11630 38528 11636
rect 38384 10804 38436 10810
rect 38384 10746 38436 10752
rect 38292 10600 38344 10606
rect 38292 10542 38344 10548
rect 38304 9994 38332 10542
rect 38108 9988 38160 9994
rect 38108 9930 38160 9936
rect 38292 9988 38344 9994
rect 38292 9930 38344 9936
rect 38120 9586 38148 9930
rect 38108 9580 38160 9586
rect 38108 9522 38160 9528
rect 38120 9450 38148 9522
rect 38198 9480 38254 9489
rect 38108 9444 38160 9450
rect 38198 9415 38200 9424
rect 38108 9386 38160 9392
rect 38252 9415 38254 9424
rect 38200 9386 38252 9392
rect 38212 8498 38240 9386
rect 38396 9178 38424 10746
rect 38488 10606 38516 11630
rect 38672 11370 38700 11698
rect 38568 11348 38620 11354
rect 38672 11342 38792 11370
rect 38568 11290 38620 11296
rect 38580 10674 38608 11290
rect 38660 11212 38712 11218
rect 38660 11154 38712 11160
rect 38568 10668 38620 10674
rect 38568 10610 38620 10616
rect 38476 10600 38528 10606
rect 38476 10542 38528 10548
rect 38488 10146 38516 10542
rect 38672 10266 38700 11154
rect 38764 10266 38792 11342
rect 38660 10260 38712 10266
rect 38660 10202 38712 10208
rect 38752 10260 38804 10266
rect 38752 10202 38804 10208
rect 38488 10118 38608 10146
rect 38580 9382 38608 10118
rect 38764 9518 38792 10202
rect 38856 10062 38884 12378
rect 38948 11626 38976 12718
rect 39132 11830 39160 13398
rect 39212 12844 39264 12850
rect 39212 12786 39264 12792
rect 39028 11824 39080 11830
rect 39028 11766 39080 11772
rect 39120 11824 39172 11830
rect 39120 11766 39172 11772
rect 38936 11620 38988 11626
rect 38936 11562 38988 11568
rect 39040 11150 39068 11766
rect 39028 11144 39080 11150
rect 39028 11086 39080 11092
rect 39132 10962 39160 11766
rect 39224 11558 39252 12786
rect 39316 12646 39344 14418
rect 39960 14414 39988 15030
rect 39948 14408 40000 14414
rect 39948 14350 40000 14356
rect 39856 13932 39908 13938
rect 39856 13874 39908 13880
rect 39868 13841 39896 13874
rect 39854 13832 39910 13841
rect 39854 13767 39910 13776
rect 40224 13728 40276 13734
rect 40224 13670 40276 13676
rect 40236 13258 40264 13670
rect 40328 13530 40356 16526
rect 40604 14618 40632 18702
rect 41156 18426 41184 19314
rect 41144 18420 41196 18426
rect 41144 18362 41196 18368
rect 41432 18290 41460 19314
rect 41800 18834 41828 19332
rect 41880 19314 41932 19320
rect 41788 18828 41840 18834
rect 41788 18770 41840 18776
rect 41800 18358 41828 18770
rect 41788 18352 41840 18358
rect 41788 18294 41840 18300
rect 41420 18284 41472 18290
rect 41420 18226 41472 18232
rect 40684 17536 40736 17542
rect 40684 17478 40736 17484
rect 40696 17270 40724 17478
rect 41144 17332 41196 17338
rect 41144 17274 41196 17280
rect 40684 17264 40736 17270
rect 40684 17206 40736 17212
rect 40868 16992 40920 16998
rect 40868 16934 40920 16940
rect 40880 16250 40908 16934
rect 41156 16250 41184 17274
rect 41432 16250 41460 18226
rect 41512 16992 41564 16998
rect 41512 16934 41564 16940
rect 41524 16590 41552 16934
rect 41512 16584 41564 16590
rect 41512 16526 41564 16532
rect 41972 16584 42024 16590
rect 41972 16526 42024 16532
rect 40868 16244 40920 16250
rect 40868 16186 40920 16192
rect 41144 16244 41196 16250
rect 41144 16186 41196 16192
rect 41420 16244 41472 16250
rect 41420 16186 41472 16192
rect 41524 16114 41552 16526
rect 41984 16114 42012 16526
rect 42076 16522 42104 21558
rect 42444 21078 42472 22170
rect 43732 21622 43760 57190
rect 49252 56710 49280 57394
rect 55508 56778 55536 57394
rect 57716 57254 57744 57394
rect 57704 57248 57756 57254
rect 57704 57190 57756 57196
rect 55496 56772 55548 56778
rect 55496 56714 55548 56720
rect 49240 56704 49292 56710
rect 49240 56646 49292 56652
rect 44824 31340 44876 31346
rect 44824 31282 44876 31288
rect 44916 31340 44968 31346
rect 44916 31282 44968 31288
rect 46756 31340 46808 31346
rect 46756 31282 46808 31288
rect 47032 31340 47084 31346
rect 47032 31282 47084 31288
rect 44836 30326 44864 31282
rect 44824 30320 44876 30326
rect 44824 30262 44876 30268
rect 44732 29708 44784 29714
rect 44732 29650 44784 29656
rect 44744 29102 44772 29650
rect 44836 29306 44864 30262
rect 44928 30122 44956 31282
rect 46296 30728 46348 30734
rect 46296 30670 46348 30676
rect 46308 30326 46336 30670
rect 46768 30394 46796 31282
rect 46940 31136 46992 31142
rect 46940 31078 46992 31084
rect 46952 30734 46980 31078
rect 46940 30728 46992 30734
rect 46940 30670 46992 30676
rect 46756 30388 46808 30394
rect 46756 30330 46808 30336
rect 46296 30320 46348 30326
rect 46296 30262 46348 30268
rect 46388 30252 46440 30258
rect 46388 30194 46440 30200
rect 44916 30116 44968 30122
rect 44916 30058 44968 30064
rect 44824 29300 44876 29306
rect 44824 29242 44876 29248
rect 44824 29164 44876 29170
rect 44824 29106 44876 29112
rect 44732 29096 44784 29102
rect 44732 29038 44784 29044
rect 44640 28076 44692 28082
rect 44640 28018 44692 28024
rect 44652 27538 44680 28018
rect 44640 27532 44692 27538
rect 44640 27474 44692 27480
rect 43904 27464 43956 27470
rect 43904 27406 43956 27412
rect 43996 27464 44048 27470
rect 43996 27406 44048 27412
rect 44180 27464 44232 27470
rect 44180 27406 44232 27412
rect 44456 27464 44508 27470
rect 44456 27406 44508 27412
rect 43916 26994 43944 27406
rect 43812 26988 43864 26994
rect 43812 26930 43864 26936
rect 43904 26988 43956 26994
rect 43904 26930 43956 26936
rect 43824 26518 43852 26930
rect 43916 26586 43944 26930
rect 43904 26580 43956 26586
rect 43904 26522 43956 26528
rect 43812 26512 43864 26518
rect 43812 26454 43864 26460
rect 43904 25832 43956 25838
rect 43904 25774 43956 25780
rect 43916 25498 43944 25774
rect 43904 25492 43956 25498
rect 43904 25434 43956 25440
rect 43812 24812 43864 24818
rect 43812 24754 43864 24760
rect 43824 24206 43852 24754
rect 43904 24608 43956 24614
rect 43904 24550 43956 24556
rect 43916 24342 43944 24550
rect 44008 24410 44036 27406
rect 44192 26858 44220 27406
rect 44468 27062 44496 27406
rect 44456 27056 44508 27062
rect 44456 26998 44508 27004
rect 44272 26920 44324 26926
rect 44272 26862 44324 26868
rect 44180 26852 44232 26858
rect 44180 26794 44232 26800
rect 44284 26314 44312 26862
rect 44468 26314 44496 26998
rect 44652 26994 44680 27474
rect 44640 26988 44692 26994
rect 44640 26930 44692 26936
rect 44272 26308 44324 26314
rect 44272 26250 44324 26256
rect 44456 26308 44508 26314
rect 44456 26250 44508 26256
rect 44284 25974 44312 26250
rect 44272 25968 44324 25974
rect 44272 25910 44324 25916
rect 44468 25362 44496 26250
rect 44744 26042 44772 29038
rect 44732 26036 44784 26042
rect 44732 25978 44784 25984
rect 44732 25900 44784 25906
rect 44732 25842 44784 25848
rect 44456 25356 44508 25362
rect 44456 25298 44508 25304
rect 44088 25152 44140 25158
rect 44088 25094 44140 25100
rect 43996 24404 44048 24410
rect 43996 24346 44048 24352
rect 43904 24336 43956 24342
rect 43904 24278 43956 24284
rect 43812 24200 43864 24206
rect 43812 24142 43864 24148
rect 43916 23866 43944 24278
rect 43904 23860 43956 23866
rect 43904 23802 43956 23808
rect 43720 21616 43772 21622
rect 43720 21558 43772 21564
rect 43444 21480 43496 21486
rect 43444 21422 43496 21428
rect 43168 21344 43220 21350
rect 43168 21286 43220 21292
rect 42432 21072 42484 21078
rect 42432 21014 42484 21020
rect 42444 20942 42472 21014
rect 42432 20936 42484 20942
rect 42432 20878 42484 20884
rect 43180 20874 43208 21286
rect 43260 21004 43312 21010
rect 43456 20992 43484 21422
rect 43312 20964 43484 20992
rect 43260 20946 43312 20952
rect 43168 20868 43220 20874
rect 43168 20810 43220 20816
rect 42616 20800 42668 20806
rect 42616 20742 42668 20748
rect 42628 20466 42656 20742
rect 42616 20460 42668 20466
rect 42616 20402 42668 20408
rect 42800 20256 42852 20262
rect 42800 20198 42852 20204
rect 42812 19922 42840 20198
rect 42800 19916 42852 19922
rect 42800 19858 42852 19864
rect 43076 19848 43128 19854
rect 43076 19790 43128 19796
rect 42248 19780 42300 19786
rect 42248 19722 42300 19728
rect 42064 16516 42116 16522
rect 42064 16458 42116 16464
rect 41512 16108 41564 16114
rect 41512 16050 41564 16056
rect 41972 16108 42024 16114
rect 41972 16050 42024 16056
rect 41604 15904 41656 15910
rect 41604 15846 41656 15852
rect 40868 15360 40920 15366
rect 40868 15302 40920 15308
rect 40592 14612 40644 14618
rect 40592 14554 40644 14560
rect 40592 14476 40644 14482
rect 40592 14418 40644 14424
rect 40500 13932 40552 13938
rect 40500 13874 40552 13880
rect 40408 13864 40460 13870
rect 40512 13841 40540 13874
rect 40408 13806 40460 13812
rect 40498 13832 40554 13841
rect 40316 13524 40368 13530
rect 40316 13466 40368 13472
rect 40420 13394 40448 13806
rect 40498 13767 40554 13776
rect 40408 13388 40460 13394
rect 40408 13330 40460 13336
rect 40224 13252 40276 13258
rect 40224 13194 40276 13200
rect 40236 12986 40264 13194
rect 40224 12980 40276 12986
rect 40224 12922 40276 12928
rect 39396 12912 39448 12918
rect 39396 12854 39448 12860
rect 39304 12640 39356 12646
rect 39304 12582 39356 12588
rect 39212 11552 39264 11558
rect 39212 11494 39264 11500
rect 39040 10934 39160 10962
rect 38936 10668 38988 10674
rect 38936 10610 38988 10616
rect 38844 10056 38896 10062
rect 38844 9998 38896 10004
rect 38752 9512 38804 9518
rect 38752 9454 38804 9460
rect 38568 9376 38620 9382
rect 38568 9318 38620 9324
rect 38384 9172 38436 9178
rect 38384 9114 38436 9120
rect 38384 8900 38436 8906
rect 38384 8842 38436 8848
rect 38200 8492 38252 8498
rect 38200 8434 38252 8440
rect 37936 7942 38056 7970
rect 37936 6497 37964 7942
rect 38016 7880 38068 7886
rect 38016 7822 38068 7828
rect 38028 7478 38056 7822
rect 38212 7750 38240 8434
rect 38396 7857 38424 8842
rect 38580 8498 38608 9318
rect 38842 9208 38898 9217
rect 38842 9143 38844 9152
rect 38896 9143 38898 9152
rect 38844 9114 38896 9120
rect 38948 9058 38976 10610
rect 38856 9030 38976 9058
rect 38568 8492 38620 8498
rect 38568 8434 38620 8440
rect 38660 8424 38712 8430
rect 38660 8366 38712 8372
rect 38672 8090 38700 8366
rect 38856 8294 38884 9030
rect 38936 8968 38988 8974
rect 38936 8910 38988 8916
rect 38948 8634 38976 8910
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 38844 8288 38896 8294
rect 38844 8230 38896 8236
rect 39040 8090 39068 10934
rect 39224 10062 39252 11494
rect 39316 10606 39344 12582
rect 39408 12442 39436 12854
rect 40132 12708 40184 12714
rect 40132 12650 40184 12656
rect 40040 12640 40092 12646
rect 40040 12582 40092 12588
rect 39396 12436 39448 12442
rect 39396 12378 39448 12384
rect 40052 12374 40080 12582
rect 40040 12368 40092 12374
rect 40040 12310 40092 12316
rect 40144 12238 40172 12650
rect 40132 12232 40184 12238
rect 40132 12174 40184 12180
rect 40236 11898 40264 12922
rect 40420 12714 40448 13330
rect 40512 12986 40540 13767
rect 40500 12980 40552 12986
rect 40500 12922 40552 12928
rect 40408 12708 40460 12714
rect 40408 12650 40460 12656
rect 40406 12336 40462 12345
rect 40406 12271 40462 12280
rect 40420 12238 40448 12271
rect 40316 12232 40368 12238
rect 40316 12174 40368 12180
rect 40408 12232 40460 12238
rect 40408 12174 40460 12180
rect 40224 11892 40276 11898
rect 40224 11834 40276 11840
rect 40328 11830 40356 12174
rect 40512 12050 40540 12922
rect 40604 12442 40632 14418
rect 40776 13184 40828 13190
rect 40776 13126 40828 13132
rect 40684 12776 40736 12782
rect 40684 12718 40736 12724
rect 40592 12436 40644 12442
rect 40592 12378 40644 12384
rect 40696 12374 40724 12718
rect 40684 12368 40736 12374
rect 40684 12310 40736 12316
rect 40420 12022 40540 12050
rect 40316 11824 40368 11830
rect 40316 11766 40368 11772
rect 40132 11756 40184 11762
rect 40132 11698 40184 11704
rect 39396 11280 39448 11286
rect 39396 11222 39448 11228
rect 39408 10674 39436 11222
rect 40144 11064 40172 11698
rect 40420 11642 40448 12022
rect 40500 11892 40552 11898
rect 40500 11834 40552 11840
rect 40328 11614 40448 11642
rect 40224 11076 40276 11082
rect 40144 11036 40224 11064
rect 40224 11018 40276 11024
rect 40236 10810 40264 11018
rect 40224 10804 40276 10810
rect 40224 10746 40276 10752
rect 39396 10668 39448 10674
rect 39396 10610 39448 10616
rect 39304 10600 39356 10606
rect 39304 10542 39356 10548
rect 39120 10056 39172 10062
rect 39120 9998 39172 10004
rect 39212 10056 39264 10062
rect 39212 9998 39264 10004
rect 38660 8084 38712 8090
rect 38660 8026 38712 8032
rect 39028 8084 39080 8090
rect 39028 8026 39080 8032
rect 38936 8016 38988 8022
rect 38936 7958 38988 7964
rect 38382 7848 38438 7857
rect 38382 7783 38438 7792
rect 38200 7744 38252 7750
rect 38200 7686 38252 7692
rect 38948 7546 38976 7958
rect 38936 7540 38988 7546
rect 38936 7482 38988 7488
rect 38016 7472 38068 7478
rect 38016 7414 38068 7420
rect 38028 7342 38056 7414
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 38660 7404 38712 7410
rect 38660 7346 38712 7352
rect 38016 7336 38068 7342
rect 38016 7278 38068 7284
rect 38028 6798 38056 7278
rect 38304 6934 38332 7346
rect 38568 7200 38620 7206
rect 38568 7142 38620 7148
rect 38292 6928 38344 6934
rect 38292 6870 38344 6876
rect 38016 6792 38068 6798
rect 38016 6734 38068 6740
rect 37922 6488 37978 6497
rect 37922 6423 37978 6432
rect 37936 6254 37964 6423
rect 38028 6390 38056 6734
rect 38016 6384 38068 6390
rect 38016 6326 38068 6332
rect 38200 6384 38252 6390
rect 38200 6326 38252 6332
rect 38108 6316 38160 6322
rect 38108 6258 38160 6264
rect 37924 6248 37976 6254
rect 37924 6190 37976 6196
rect 38016 6112 38068 6118
rect 37844 6072 37964 6100
rect 37830 5536 37886 5545
rect 37830 5471 37886 5480
rect 37844 4826 37872 5471
rect 37936 5234 37964 6072
rect 38016 6054 38068 6060
rect 38028 5710 38056 6054
rect 38016 5704 38068 5710
rect 38016 5646 38068 5652
rect 38014 5400 38070 5409
rect 38014 5335 38070 5344
rect 37924 5228 37976 5234
rect 37924 5170 37976 5176
rect 38028 5166 38056 5335
rect 38016 5160 38068 5166
rect 38016 5102 38068 5108
rect 37832 4820 37884 4826
rect 37832 4762 37884 4768
rect 38120 4622 38148 6258
rect 38212 5710 38240 6326
rect 38304 6118 38332 6870
rect 38580 6202 38608 7142
rect 38672 7002 38700 7346
rect 38660 6996 38712 7002
rect 38660 6938 38712 6944
rect 39132 6662 39160 9998
rect 39408 9654 39436 10610
rect 39764 10600 39816 10606
rect 39764 10542 39816 10548
rect 39776 9722 39804 10542
rect 40224 10056 40276 10062
rect 40224 9998 40276 10004
rect 39764 9716 39816 9722
rect 39764 9658 39816 9664
rect 39396 9648 39448 9654
rect 39396 9590 39448 9596
rect 39580 9580 39632 9586
rect 39580 9522 39632 9528
rect 39592 9042 39620 9522
rect 39580 9036 39632 9042
rect 39580 8978 39632 8984
rect 39776 8906 39804 9658
rect 40236 9586 40264 9998
rect 40224 9580 40276 9586
rect 40224 9522 40276 9528
rect 39764 8900 39816 8906
rect 39764 8842 39816 8848
rect 40132 8832 40184 8838
rect 40132 8774 40184 8780
rect 39396 8492 39448 8498
rect 39396 8434 39448 8440
rect 39580 8492 39632 8498
rect 39580 8434 39632 8440
rect 39408 8022 39436 8434
rect 39396 8016 39448 8022
rect 39396 7958 39448 7964
rect 39592 7954 39620 8434
rect 39580 7948 39632 7954
rect 39580 7890 39632 7896
rect 39592 7478 39620 7890
rect 39580 7472 39632 7478
rect 39580 7414 39632 7420
rect 39396 7336 39448 7342
rect 39396 7278 39448 7284
rect 39120 6656 39172 6662
rect 39120 6598 39172 6604
rect 39304 6656 39356 6662
rect 39304 6598 39356 6604
rect 38660 6384 38712 6390
rect 38658 6352 38660 6361
rect 38844 6384 38896 6390
rect 38712 6352 38714 6361
rect 38844 6326 38896 6332
rect 38658 6287 38714 6296
rect 38580 6186 38700 6202
rect 38856 6186 38884 6326
rect 38936 6316 38988 6322
rect 38936 6258 38988 6264
rect 39120 6316 39172 6322
rect 39120 6258 39172 6264
rect 38580 6180 38712 6186
rect 38580 6174 38660 6180
rect 38660 6122 38712 6128
rect 38844 6180 38896 6186
rect 38844 6122 38896 6128
rect 38292 6112 38344 6118
rect 38292 6054 38344 6060
rect 38290 5808 38346 5817
rect 38290 5743 38346 5752
rect 38304 5710 38332 5743
rect 38200 5704 38252 5710
rect 38200 5646 38252 5652
rect 38292 5704 38344 5710
rect 38292 5646 38344 5652
rect 38476 5704 38528 5710
rect 38476 5646 38528 5652
rect 38212 5302 38240 5646
rect 38200 5296 38252 5302
rect 38200 5238 38252 5244
rect 38108 4616 38160 4622
rect 38108 4558 38160 4564
rect 37740 4072 37792 4078
rect 37740 4014 37792 4020
rect 38304 3942 38332 5646
rect 38488 5234 38516 5646
rect 38476 5228 38528 5234
rect 38476 5170 38528 5176
rect 38568 5160 38620 5166
rect 38568 5102 38620 5108
rect 38580 4758 38608 5102
rect 38948 5098 38976 6258
rect 39132 5710 39160 6258
rect 39120 5704 39172 5710
rect 39120 5646 39172 5652
rect 38936 5092 38988 5098
rect 38936 5034 38988 5040
rect 38568 4752 38620 4758
rect 38568 4694 38620 4700
rect 38476 4072 38528 4078
rect 38476 4014 38528 4020
rect 38292 3936 38344 3942
rect 38292 3878 38344 3884
rect 37648 3188 37700 3194
rect 37648 3130 37700 3136
rect 38488 3058 38516 4014
rect 38476 3052 38528 3058
rect 38476 2994 38528 3000
rect 37556 2984 37608 2990
rect 37556 2926 37608 2932
rect 38108 2984 38160 2990
rect 38108 2926 38160 2932
rect 36096 2746 36308 2774
rect 37292 2746 37504 2774
rect 36280 2650 36308 2746
rect 36268 2644 36320 2650
rect 36268 2586 36320 2592
rect 37476 2514 37504 2746
rect 38120 2650 38148 2926
rect 38108 2644 38160 2650
rect 38108 2586 38160 2592
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 34428 2304 34480 2310
rect 34428 2246 34480 2252
rect 38580 2038 38608 4694
rect 39316 3126 39344 6598
rect 39408 5710 39436 7278
rect 39488 6792 39540 6798
rect 39488 6734 39540 6740
rect 39500 5914 39528 6734
rect 39856 6452 39908 6458
rect 39856 6394 39908 6400
rect 39868 6322 39896 6394
rect 39856 6316 39908 6322
rect 39856 6258 39908 6264
rect 39868 6118 39896 6258
rect 39856 6112 39908 6118
rect 39856 6054 39908 6060
rect 39488 5908 39540 5914
rect 39488 5850 39540 5856
rect 39396 5704 39448 5710
rect 39396 5646 39448 5652
rect 40040 5704 40092 5710
rect 40040 5646 40092 5652
rect 40052 5302 40080 5646
rect 40040 5296 40092 5302
rect 40040 5238 40092 5244
rect 40052 4214 40080 5238
rect 40040 4208 40092 4214
rect 40040 4150 40092 4156
rect 40040 4072 40092 4078
rect 40040 4014 40092 4020
rect 40052 3738 40080 4014
rect 40040 3732 40092 3738
rect 40040 3674 40092 3680
rect 40144 3398 40172 8774
rect 40224 8016 40276 8022
rect 40224 7958 40276 7964
rect 40236 6798 40264 7958
rect 40224 6792 40276 6798
rect 40224 6734 40276 6740
rect 40236 4690 40264 6734
rect 40224 4684 40276 4690
rect 40224 4626 40276 4632
rect 40328 4298 40356 11614
rect 40408 11552 40460 11558
rect 40408 11494 40460 11500
rect 40420 11150 40448 11494
rect 40408 11144 40460 11150
rect 40408 11086 40460 11092
rect 40408 9988 40460 9994
rect 40408 9930 40460 9936
rect 40420 9042 40448 9930
rect 40408 9036 40460 9042
rect 40408 8978 40460 8984
rect 40408 8900 40460 8906
rect 40408 8842 40460 8848
rect 40420 8294 40448 8842
rect 40408 8288 40460 8294
rect 40408 8230 40460 8236
rect 40420 7546 40448 8230
rect 40512 8090 40540 11834
rect 40788 11354 40816 13126
rect 40776 11348 40828 11354
rect 40776 11290 40828 11296
rect 40684 10668 40736 10674
rect 40684 10610 40736 10616
rect 40696 9178 40724 10610
rect 40684 9172 40736 9178
rect 40684 9114 40736 9120
rect 40592 9104 40644 9110
rect 40592 9046 40644 9052
rect 40604 8498 40632 9046
rect 40592 8492 40644 8498
rect 40592 8434 40644 8440
rect 40500 8084 40552 8090
rect 40500 8026 40552 8032
rect 40408 7540 40460 7546
rect 40408 7482 40460 7488
rect 40512 7274 40540 8026
rect 40696 7478 40724 9114
rect 40776 8356 40828 8362
rect 40776 8298 40828 8304
rect 40684 7472 40736 7478
rect 40684 7414 40736 7420
rect 40696 7274 40724 7414
rect 40500 7268 40552 7274
rect 40500 7210 40552 7216
rect 40684 7268 40736 7274
rect 40684 7210 40736 7216
rect 40512 6798 40540 7210
rect 40500 6792 40552 6798
rect 40500 6734 40552 6740
rect 40408 6656 40460 6662
rect 40408 6598 40460 6604
rect 40420 6361 40448 6598
rect 40406 6352 40462 6361
rect 40406 6287 40408 6296
rect 40460 6287 40462 6296
rect 40408 6258 40460 6264
rect 40420 6227 40448 6258
rect 40684 5840 40736 5846
rect 40684 5782 40736 5788
rect 40696 5574 40724 5782
rect 40684 5568 40736 5574
rect 40684 5510 40736 5516
rect 40592 5160 40644 5166
rect 40592 5102 40644 5108
rect 40500 5024 40552 5030
rect 40500 4966 40552 4972
rect 40236 4270 40356 4298
rect 40132 3392 40184 3398
rect 40132 3334 40184 3340
rect 39304 3120 39356 3126
rect 39304 3062 39356 3068
rect 40236 2990 40264 4270
rect 40316 4208 40368 4214
rect 40368 4168 40448 4196
rect 40316 4150 40368 4156
rect 40316 3528 40368 3534
rect 40316 3470 40368 3476
rect 40328 3194 40356 3470
rect 40316 3188 40368 3194
rect 40316 3130 40368 3136
rect 40420 3126 40448 4168
rect 40512 3534 40540 4966
rect 40604 3602 40632 5102
rect 40696 4978 40724 5510
rect 40788 5098 40816 8298
rect 40776 5092 40828 5098
rect 40776 5034 40828 5040
rect 40696 4950 40816 4978
rect 40684 4480 40736 4486
rect 40684 4422 40736 4428
rect 40592 3596 40644 3602
rect 40592 3538 40644 3544
rect 40500 3528 40552 3534
rect 40500 3470 40552 3476
rect 40604 3126 40632 3538
rect 40408 3120 40460 3126
rect 40408 3062 40460 3068
rect 40592 3120 40644 3126
rect 40592 3062 40644 3068
rect 40224 2984 40276 2990
rect 40224 2926 40276 2932
rect 40040 2848 40092 2854
rect 40040 2790 40092 2796
rect 40052 2446 40080 2790
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 40696 2378 40724 4422
rect 40788 2990 40816 4950
rect 40880 4282 40908 15302
rect 41420 15088 41472 15094
rect 41420 15030 41472 15036
rect 41432 14618 41460 15030
rect 41420 14612 41472 14618
rect 41420 14554 41472 14560
rect 41616 14074 41644 15846
rect 41984 15162 42012 16050
rect 41972 15156 42024 15162
rect 41972 15098 42024 15104
rect 41696 14408 41748 14414
rect 41696 14350 41748 14356
rect 41604 14068 41656 14074
rect 41604 14010 41656 14016
rect 41708 13870 41736 14350
rect 41972 14272 42024 14278
rect 41972 14214 42024 14220
rect 41696 13864 41748 13870
rect 41696 13806 41748 13812
rect 41236 13388 41288 13394
rect 41236 13330 41288 13336
rect 41248 12102 41276 13330
rect 41984 13326 42012 14214
rect 41972 13320 42024 13326
rect 41972 13262 42024 13268
rect 41984 12782 42012 13262
rect 41972 12776 42024 12782
rect 41972 12718 42024 12724
rect 40960 12096 41012 12102
rect 40960 12038 41012 12044
rect 41236 12096 41288 12102
rect 41236 12038 41288 12044
rect 40972 9450 41000 12038
rect 41248 10130 41276 12038
rect 41788 11008 41840 11014
rect 41788 10950 41840 10956
rect 41800 10742 41828 10950
rect 41788 10736 41840 10742
rect 41788 10678 41840 10684
rect 41236 10124 41288 10130
rect 41236 10066 41288 10072
rect 41248 9586 41276 10066
rect 41328 10056 41380 10062
rect 41326 10024 41328 10033
rect 41380 10024 41382 10033
rect 41326 9959 41382 9968
rect 41326 9616 41382 9625
rect 41236 9580 41288 9586
rect 41326 9551 41382 9560
rect 41236 9522 41288 9528
rect 40960 9444 41012 9450
rect 40960 9386 41012 9392
rect 40972 8090 41000 9386
rect 41340 9042 41368 9551
rect 41328 9036 41380 9042
rect 41328 8978 41380 8984
rect 41052 8968 41104 8974
rect 41052 8910 41104 8916
rect 41144 8968 41196 8974
rect 41144 8910 41196 8916
rect 40960 8084 41012 8090
rect 40960 8026 41012 8032
rect 40960 7404 41012 7410
rect 40960 7346 41012 7352
rect 40972 6458 41000 7346
rect 41064 7206 41092 8910
rect 41052 7200 41104 7206
rect 41052 7142 41104 7148
rect 41156 7002 41184 8910
rect 41340 8090 41368 8978
rect 41788 8968 41840 8974
rect 41788 8910 41840 8916
rect 42156 8968 42208 8974
rect 42156 8910 42208 8916
rect 41800 8498 41828 8910
rect 42168 8498 42196 8910
rect 41788 8492 41840 8498
rect 41788 8434 41840 8440
rect 42156 8492 42208 8498
rect 42156 8434 42208 8440
rect 41604 8356 41656 8362
rect 41604 8298 41656 8304
rect 41328 8084 41380 8090
rect 41328 8026 41380 8032
rect 41420 7880 41472 7886
rect 41420 7822 41472 7828
rect 41144 6996 41196 7002
rect 41064 6956 41144 6984
rect 40960 6452 41012 6458
rect 40960 6394 41012 6400
rect 41064 6322 41092 6956
rect 41144 6938 41196 6944
rect 41432 6798 41460 7822
rect 41616 7818 41644 8298
rect 42156 7948 42208 7954
rect 42156 7890 42208 7896
rect 41604 7812 41656 7818
rect 41604 7754 41656 7760
rect 41512 7744 41564 7750
rect 41512 7686 41564 7692
rect 41420 6792 41472 6798
rect 41420 6734 41472 6740
rect 41432 6662 41460 6734
rect 41420 6656 41472 6662
rect 41420 6598 41472 6604
rect 41052 6316 41104 6322
rect 40972 6276 41052 6304
rect 40972 5166 41000 6276
rect 41052 6258 41104 6264
rect 41144 6248 41196 6254
rect 41144 6190 41196 6196
rect 41156 5710 41184 6190
rect 41432 5846 41460 6598
rect 41524 6458 41552 7686
rect 41616 6934 41644 7754
rect 41972 7200 42024 7206
rect 41972 7142 42024 7148
rect 41604 6928 41656 6934
rect 41604 6870 41656 6876
rect 41984 6866 42012 7142
rect 41972 6860 42024 6866
rect 41972 6802 42024 6808
rect 41512 6452 41564 6458
rect 41512 6394 41564 6400
rect 41420 5840 41472 5846
rect 41420 5782 41472 5788
rect 41144 5704 41196 5710
rect 41144 5646 41196 5652
rect 41328 5704 41380 5710
rect 41328 5646 41380 5652
rect 41052 5568 41104 5574
rect 41052 5510 41104 5516
rect 41064 5302 41092 5510
rect 41052 5296 41104 5302
rect 41052 5238 41104 5244
rect 40960 5160 41012 5166
rect 40960 5102 41012 5108
rect 40868 4276 40920 4282
rect 40868 4218 40920 4224
rect 40880 3058 40908 4218
rect 40868 3052 40920 3058
rect 40868 2994 40920 3000
rect 40972 2990 41000 5102
rect 41156 4146 41184 5646
rect 41236 5636 41288 5642
rect 41236 5578 41288 5584
rect 41144 4140 41196 4146
rect 41144 4082 41196 4088
rect 41248 3602 41276 5578
rect 41340 4826 41368 5646
rect 41418 5264 41474 5273
rect 41418 5199 41420 5208
rect 41472 5199 41474 5208
rect 41420 5170 41472 5176
rect 41328 4820 41380 4826
rect 41328 4762 41380 4768
rect 41524 4486 41552 6394
rect 42168 5914 42196 7890
rect 42156 5908 42208 5914
rect 42156 5850 42208 5856
rect 42064 5636 42116 5642
rect 42064 5578 42116 5584
rect 41788 5296 41840 5302
rect 41788 5238 41840 5244
rect 41604 5160 41656 5166
rect 41604 5102 41656 5108
rect 41616 5030 41644 5102
rect 41604 5024 41656 5030
rect 41604 4966 41656 4972
rect 41696 4684 41748 4690
rect 41696 4626 41748 4632
rect 41512 4480 41564 4486
rect 41512 4422 41564 4428
rect 41524 4162 41552 4422
rect 41708 4214 41736 4626
rect 41432 4134 41552 4162
rect 41696 4208 41748 4214
rect 41696 4150 41748 4156
rect 41432 4026 41460 4134
rect 41340 3998 41460 4026
rect 41510 4040 41566 4049
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 40776 2984 40828 2990
rect 40776 2926 40828 2932
rect 40960 2984 41012 2990
rect 40960 2926 41012 2932
rect 41340 2650 41368 3998
rect 41510 3975 41512 3984
rect 41564 3975 41566 3984
rect 41512 3946 41564 3952
rect 41800 3194 41828 5238
rect 42076 5166 42104 5578
rect 42064 5160 42116 5166
rect 42064 5102 42116 5108
rect 41880 4820 41932 4826
rect 41880 4762 41932 4768
rect 41892 4622 41920 4762
rect 42076 4622 42104 5102
rect 42154 4720 42210 4729
rect 42154 4655 42156 4664
rect 42208 4655 42210 4664
rect 42156 4626 42208 4632
rect 41880 4616 41932 4622
rect 41880 4558 41932 4564
rect 42064 4616 42116 4622
rect 42064 4558 42116 4564
rect 41788 3188 41840 3194
rect 41788 3130 41840 3136
rect 41328 2644 41380 2650
rect 41328 2586 41380 2592
rect 42260 2514 42288 19722
rect 43088 19514 43116 19790
rect 43076 19508 43128 19514
rect 43076 19450 43128 19456
rect 42800 19372 42852 19378
rect 42800 19314 42852 19320
rect 42812 18970 42840 19314
rect 42800 18964 42852 18970
rect 42800 18906 42852 18912
rect 43180 18630 43208 20810
rect 43456 20602 43484 20964
rect 43444 20596 43496 20602
rect 43444 20538 43496 20544
rect 43720 19712 43772 19718
rect 43720 19654 43772 19660
rect 43732 19514 43760 19654
rect 43720 19508 43772 19514
rect 43720 19450 43772 19456
rect 43626 19408 43682 19417
rect 44100 19378 44128 25094
rect 44272 24676 44324 24682
rect 44272 24618 44324 24624
rect 44180 24132 44232 24138
rect 44180 24074 44232 24080
rect 44192 23730 44220 24074
rect 44180 23724 44232 23730
rect 44180 23666 44232 23672
rect 44192 22778 44220 23666
rect 44284 23118 44312 24618
rect 44468 23730 44496 25298
rect 44744 24614 44772 25842
rect 44732 24608 44784 24614
rect 44732 24550 44784 24556
rect 44456 23724 44508 23730
rect 44456 23666 44508 23672
rect 44468 23526 44496 23666
rect 44456 23520 44508 23526
rect 44456 23462 44508 23468
rect 44364 23180 44416 23186
rect 44364 23122 44416 23128
rect 44272 23112 44324 23118
rect 44272 23054 44324 23060
rect 44180 22772 44232 22778
rect 44180 22714 44232 22720
rect 43626 19343 43628 19352
rect 43680 19343 43682 19352
rect 44088 19372 44140 19378
rect 43628 19314 43680 19320
rect 44088 19314 44140 19320
rect 43996 19304 44048 19310
rect 43996 19246 44048 19252
rect 43260 19168 43312 19174
rect 43260 19110 43312 19116
rect 43272 18766 43300 19110
rect 43260 18760 43312 18766
rect 43260 18702 43312 18708
rect 44008 18630 44036 19246
rect 43168 18624 43220 18630
rect 43168 18566 43220 18572
rect 43996 18624 44048 18630
rect 43996 18566 44048 18572
rect 43720 18284 43772 18290
rect 43720 18226 43772 18232
rect 43732 17678 43760 18226
rect 43904 18080 43956 18086
rect 43902 18048 43904 18057
rect 43956 18048 43958 18057
rect 43902 17983 43958 17992
rect 43444 17672 43496 17678
rect 43444 17614 43496 17620
rect 43720 17672 43772 17678
rect 43720 17614 43772 17620
rect 42708 17536 42760 17542
rect 42708 17478 42760 17484
rect 42720 17202 42748 17478
rect 43456 17338 43484 17614
rect 43536 17604 43588 17610
rect 43536 17546 43588 17552
rect 43548 17338 43576 17546
rect 43444 17332 43496 17338
rect 43444 17274 43496 17280
rect 43536 17332 43588 17338
rect 43536 17274 43588 17280
rect 42708 17196 42760 17202
rect 42708 17138 42760 17144
rect 43444 17196 43496 17202
rect 43444 17138 43496 17144
rect 42524 16992 42576 16998
rect 42524 16934 42576 16940
rect 42536 16046 42564 16934
rect 42720 16794 42748 17138
rect 42708 16788 42760 16794
rect 42708 16730 42760 16736
rect 42800 16244 42852 16250
rect 42800 16186 42852 16192
rect 42708 16108 42760 16114
rect 42708 16050 42760 16056
rect 42524 16040 42576 16046
rect 42524 15982 42576 15988
rect 42536 15434 42564 15982
rect 42524 15428 42576 15434
rect 42524 15370 42576 15376
rect 42536 14414 42564 15370
rect 42524 14408 42576 14414
rect 42524 14350 42576 14356
rect 42340 13864 42392 13870
rect 42340 13806 42392 13812
rect 42352 13190 42380 13806
rect 42340 13184 42392 13190
rect 42340 13126 42392 13132
rect 42340 11756 42392 11762
rect 42340 11698 42392 11704
rect 42352 11354 42380 11698
rect 42340 11348 42392 11354
rect 42340 11290 42392 11296
rect 42352 10742 42380 11290
rect 42340 10736 42392 10742
rect 42340 10678 42392 10684
rect 42432 10668 42484 10674
rect 42432 10610 42484 10616
rect 42444 9382 42472 10610
rect 42432 9376 42484 9382
rect 42432 9318 42484 9324
rect 42536 9110 42564 14350
rect 42720 12986 42748 16050
rect 42812 15638 42840 16186
rect 42800 15632 42852 15638
rect 42800 15574 42852 15580
rect 43260 15496 43312 15502
rect 43260 15438 43312 15444
rect 43076 14612 43128 14618
rect 43076 14554 43128 14560
rect 42984 14000 43036 14006
rect 42984 13942 43036 13948
rect 42996 13326 43024 13942
rect 43088 13530 43116 14554
rect 43272 14550 43300 15438
rect 43456 15162 43484 17138
rect 43626 16008 43682 16017
rect 43626 15943 43628 15952
rect 43680 15943 43682 15952
rect 43628 15914 43680 15920
rect 43628 15428 43680 15434
rect 43628 15370 43680 15376
rect 43444 15156 43496 15162
rect 43444 15098 43496 15104
rect 43536 15020 43588 15026
rect 43536 14962 43588 14968
rect 43640 15008 43668 15370
rect 43732 15162 43760 17614
rect 43812 17196 43864 17202
rect 43812 17138 43864 17144
rect 43824 16522 43852 17138
rect 43812 16516 43864 16522
rect 43812 16458 43864 16464
rect 43824 16250 43852 16458
rect 43812 16244 43864 16250
rect 43812 16186 43864 16192
rect 43720 15156 43772 15162
rect 43720 15098 43772 15104
rect 43720 15020 43772 15026
rect 43640 14980 43720 15008
rect 43260 14544 43312 14550
rect 43260 14486 43312 14492
rect 43444 14272 43496 14278
rect 43548 14260 43576 14962
rect 43496 14232 43576 14260
rect 43444 14214 43496 14220
rect 43548 14074 43576 14232
rect 43536 14068 43588 14074
rect 43536 14010 43588 14016
rect 43640 13954 43668 14980
rect 43720 14962 43772 14968
rect 43824 14822 43852 16186
rect 43904 14884 43956 14890
rect 43904 14826 43956 14832
rect 43812 14816 43864 14822
rect 43812 14758 43864 14764
rect 43824 13954 43852 14758
rect 43916 14414 43944 14826
rect 43904 14408 43956 14414
rect 43904 14350 43956 14356
rect 43352 13932 43404 13938
rect 43352 13874 43404 13880
rect 43456 13926 43668 13954
rect 43732 13926 43852 13954
rect 43076 13524 43128 13530
rect 43076 13466 43128 13472
rect 43364 13394 43392 13874
rect 43352 13388 43404 13394
rect 43352 13330 43404 13336
rect 42984 13320 43036 13326
rect 42890 13288 42946 13297
rect 42984 13262 43036 13268
rect 43168 13320 43220 13326
rect 43168 13262 43220 13268
rect 42890 13223 42946 13232
rect 42708 12980 42760 12986
rect 42708 12922 42760 12928
rect 42616 12912 42668 12918
rect 42616 12854 42668 12860
rect 42628 11150 42656 12854
rect 42904 12850 42932 13223
rect 42892 12844 42944 12850
rect 42892 12786 42944 12792
rect 42996 12434 43024 13262
rect 43076 12844 43128 12850
rect 43076 12786 43128 12792
rect 42904 12406 43024 12434
rect 42800 11688 42852 11694
rect 42800 11630 42852 11636
rect 42708 11212 42760 11218
rect 42708 11154 42760 11160
rect 42616 11144 42668 11150
rect 42616 11086 42668 11092
rect 42616 9376 42668 9382
rect 42616 9318 42668 9324
rect 42524 9104 42576 9110
rect 42524 9046 42576 9052
rect 42524 8084 42576 8090
rect 42524 8026 42576 8032
rect 42536 7342 42564 8026
rect 42524 7336 42576 7342
rect 42524 7278 42576 7284
rect 42536 6866 42564 7278
rect 42524 6860 42576 6866
rect 42524 6802 42576 6808
rect 42524 6316 42576 6322
rect 42524 6258 42576 6264
rect 42340 5568 42392 5574
rect 42340 5510 42392 5516
rect 42352 4554 42380 5510
rect 42432 4820 42484 4826
rect 42432 4762 42484 4768
rect 42444 4690 42472 4762
rect 42536 4758 42564 6258
rect 42628 6202 42656 9318
rect 42720 7954 42748 11154
rect 42812 9110 42840 11630
rect 42800 9104 42852 9110
rect 42800 9046 42852 9052
rect 42800 8016 42852 8022
rect 42800 7958 42852 7964
rect 42708 7948 42760 7954
rect 42708 7890 42760 7896
rect 42812 7546 42840 7958
rect 42800 7540 42852 7546
rect 42800 7482 42852 7488
rect 42904 7410 42932 12406
rect 43088 12288 43116 12786
rect 43180 12374 43208 13262
rect 43260 12844 43312 12850
rect 43260 12786 43312 12792
rect 43168 12368 43220 12374
rect 43168 12310 43220 12316
rect 42996 12260 43116 12288
rect 42996 11762 43024 12260
rect 43168 12232 43220 12238
rect 43168 12174 43220 12180
rect 43076 12164 43128 12170
rect 43076 12106 43128 12112
rect 43088 11762 43116 12106
rect 42984 11756 43036 11762
rect 42984 11698 43036 11704
rect 43076 11756 43128 11762
rect 43076 11698 43128 11704
rect 42996 8566 43024 11698
rect 43088 11064 43116 11698
rect 43180 11218 43208 12174
rect 43272 12102 43300 12786
rect 43364 12238 43392 13330
rect 43352 12232 43404 12238
rect 43352 12174 43404 12180
rect 43260 12096 43312 12102
rect 43260 12038 43312 12044
rect 43272 11898 43300 12038
rect 43260 11892 43312 11898
rect 43260 11834 43312 11840
rect 43364 11642 43392 12174
rect 43456 11762 43484 13926
rect 43536 13796 43588 13802
rect 43536 13738 43588 13744
rect 43548 12306 43576 13738
rect 43732 13161 43760 13926
rect 43916 13394 43944 14350
rect 43904 13388 43956 13394
rect 43904 13330 43956 13336
rect 43812 13320 43864 13326
rect 43810 13288 43812 13297
rect 43864 13288 43866 13297
rect 43810 13223 43866 13232
rect 43718 13152 43774 13161
rect 43718 13087 43774 13096
rect 43916 12918 43944 13330
rect 43904 12912 43956 12918
rect 43904 12854 43956 12860
rect 43628 12844 43680 12850
rect 43628 12786 43680 12792
rect 43536 12300 43588 12306
rect 43536 12242 43588 12248
rect 43640 11830 43668 12786
rect 44008 12764 44036 18566
rect 44284 18426 44312 23054
rect 44376 22234 44404 23122
rect 44640 23112 44692 23118
rect 44640 23054 44692 23060
rect 44548 22976 44600 22982
rect 44548 22918 44600 22924
rect 44560 22234 44588 22918
rect 44364 22228 44416 22234
rect 44364 22170 44416 22176
rect 44548 22228 44600 22234
rect 44548 22170 44600 22176
rect 44456 21956 44508 21962
rect 44456 21898 44508 21904
rect 44468 21622 44496 21898
rect 44456 21616 44508 21622
rect 44456 21558 44508 21564
rect 44468 20466 44496 21558
rect 44548 20800 44600 20806
rect 44548 20742 44600 20748
rect 44456 20460 44508 20466
rect 44456 20402 44508 20408
rect 44364 20392 44416 20398
rect 44468 20369 44496 20402
rect 44364 20334 44416 20340
rect 44454 20360 44510 20369
rect 44376 20058 44404 20334
rect 44454 20295 44510 20304
rect 44364 20052 44416 20058
rect 44364 19994 44416 20000
rect 44560 19854 44588 20742
rect 44548 19848 44600 19854
rect 44548 19790 44600 19796
rect 44560 19310 44588 19790
rect 44548 19304 44600 19310
rect 44548 19246 44600 19252
rect 44272 18420 44324 18426
rect 44272 18362 44324 18368
rect 44456 18284 44508 18290
rect 44456 18226 44508 18232
rect 44180 17672 44232 17678
rect 44180 17614 44232 17620
rect 44088 16040 44140 16046
rect 44088 15982 44140 15988
rect 43824 12736 44036 12764
rect 43720 12640 43772 12646
rect 43718 12608 43720 12617
rect 43772 12608 43774 12617
rect 43718 12543 43774 12552
rect 43720 12368 43772 12374
rect 43720 12310 43772 12316
rect 43628 11824 43680 11830
rect 43628 11766 43680 11772
rect 43444 11756 43496 11762
rect 43444 11698 43496 11704
rect 43364 11614 43484 11642
rect 43352 11552 43404 11558
rect 43352 11494 43404 11500
rect 43364 11354 43392 11494
rect 43352 11348 43404 11354
rect 43352 11290 43404 11296
rect 43168 11212 43220 11218
rect 43168 11154 43220 11160
rect 43168 11076 43220 11082
rect 43088 11036 43168 11064
rect 43168 11018 43220 11024
rect 43456 10742 43484 11614
rect 43444 10736 43496 10742
rect 43444 10678 43496 10684
rect 43076 10464 43128 10470
rect 43076 10406 43128 10412
rect 42984 8560 43036 8566
rect 42984 8502 43036 8508
rect 42984 8424 43036 8430
rect 43088 8412 43116 10406
rect 43168 9988 43220 9994
rect 43168 9930 43220 9936
rect 43352 9988 43404 9994
rect 43352 9930 43404 9936
rect 43180 8838 43208 9930
rect 43364 9761 43392 9930
rect 43456 9926 43484 10678
rect 43444 9920 43496 9926
rect 43444 9862 43496 9868
rect 43350 9752 43406 9761
rect 43350 9687 43406 9696
rect 43456 8906 43484 9862
rect 43536 9104 43588 9110
rect 43536 9046 43588 9052
rect 43444 8900 43496 8906
rect 43444 8842 43496 8848
rect 43168 8832 43220 8838
rect 43168 8774 43220 8780
rect 43180 8430 43208 8774
rect 43036 8384 43116 8412
rect 43168 8424 43220 8430
rect 42984 8366 43036 8372
rect 43168 8366 43220 8372
rect 42996 7410 43024 8366
rect 43260 7744 43312 7750
rect 43260 7686 43312 7692
rect 42892 7404 42944 7410
rect 42892 7346 42944 7352
rect 42984 7404 43036 7410
rect 42984 7346 43036 7352
rect 43168 7404 43220 7410
rect 43168 7346 43220 7352
rect 42904 6866 42932 7346
rect 42892 6860 42944 6866
rect 42944 6820 43024 6848
rect 42892 6802 42944 6808
rect 42996 6730 43024 6820
rect 42984 6724 43036 6730
rect 42984 6666 43036 6672
rect 42628 6174 42748 6202
rect 42616 6112 42668 6118
rect 42616 6054 42668 6060
rect 42524 4752 42576 4758
rect 42524 4694 42576 4700
rect 42432 4684 42484 4690
rect 42432 4626 42484 4632
rect 42340 4548 42392 4554
rect 42340 4490 42392 4496
rect 42628 4146 42656 6054
rect 42720 4604 42748 6174
rect 42800 5908 42852 5914
rect 42800 5850 42852 5856
rect 42812 5302 42840 5850
rect 43180 5778 43208 7346
rect 43272 5817 43300 7686
rect 43352 7540 43404 7546
rect 43352 7482 43404 7488
rect 43258 5808 43314 5817
rect 43168 5772 43220 5778
rect 43364 5778 43392 7482
rect 43456 7342 43484 8842
rect 43548 8498 43576 9046
rect 43640 9042 43668 11766
rect 43732 11286 43760 12310
rect 43720 11280 43772 11286
rect 43720 11222 43772 11228
rect 43732 10470 43760 11222
rect 43720 10464 43772 10470
rect 43720 10406 43772 10412
rect 43718 9480 43774 9489
rect 43718 9415 43774 9424
rect 43732 9382 43760 9415
rect 43720 9376 43772 9382
rect 43720 9318 43772 9324
rect 43628 9036 43680 9042
rect 43628 8978 43680 8984
rect 43628 8900 43680 8906
rect 43628 8842 43680 8848
rect 43536 8492 43588 8498
rect 43536 8434 43588 8440
rect 43444 7336 43496 7342
rect 43444 7278 43496 7284
rect 43640 6934 43668 8842
rect 43718 7168 43774 7177
rect 43718 7103 43774 7112
rect 43732 7002 43760 7103
rect 43720 6996 43772 7002
rect 43720 6938 43772 6944
rect 43628 6928 43680 6934
rect 43628 6870 43680 6876
rect 43258 5743 43314 5752
rect 43352 5772 43404 5778
rect 43168 5714 43220 5720
rect 43272 5710 43300 5743
rect 43352 5714 43404 5720
rect 43260 5704 43312 5710
rect 43640 5658 43668 6870
rect 43260 5646 43312 5652
rect 42984 5636 43036 5642
rect 42984 5578 43036 5584
rect 43364 5630 43668 5658
rect 42800 5296 42852 5302
rect 42800 5238 42852 5244
rect 42892 4616 42944 4622
rect 42720 4576 42892 4604
rect 42892 4558 42944 4564
rect 42616 4140 42668 4146
rect 42616 4082 42668 4088
rect 42628 3602 42656 4082
rect 42616 3596 42668 3602
rect 42616 3538 42668 3544
rect 42904 2854 42932 4558
rect 42996 3126 43024 5578
rect 43364 4146 43392 5630
rect 43720 5296 43772 5302
rect 43720 5238 43772 5244
rect 43628 4752 43680 4758
rect 43628 4694 43680 4700
rect 43444 4548 43496 4554
rect 43444 4490 43496 4496
rect 43536 4548 43588 4554
rect 43536 4490 43588 4496
rect 43352 4140 43404 4146
rect 43352 4082 43404 4088
rect 43456 3942 43484 4490
rect 43548 4214 43576 4490
rect 43640 4282 43668 4694
rect 43628 4276 43680 4282
rect 43628 4218 43680 4224
rect 43732 4214 43760 5238
rect 43536 4208 43588 4214
rect 43536 4150 43588 4156
rect 43720 4208 43772 4214
rect 43720 4150 43772 4156
rect 43352 3936 43404 3942
rect 43352 3878 43404 3884
rect 43444 3936 43496 3942
rect 43444 3878 43496 3884
rect 43364 3738 43392 3878
rect 43352 3732 43404 3738
rect 43352 3674 43404 3680
rect 43536 3528 43588 3534
rect 43536 3470 43588 3476
rect 42984 3120 43036 3126
rect 42984 3062 43036 3068
rect 43260 2984 43312 2990
rect 43260 2926 43312 2932
rect 42892 2848 42944 2854
rect 42892 2790 42944 2796
rect 43272 2774 43300 2926
rect 43180 2746 43300 2774
rect 43180 2650 43208 2746
rect 43168 2644 43220 2650
rect 43168 2586 43220 2592
rect 43548 2582 43576 3470
rect 43732 3466 43760 4150
rect 43824 3534 43852 12736
rect 43994 12608 44050 12617
rect 43994 12543 44050 12552
rect 44008 12170 44036 12543
rect 44100 12442 44128 15982
rect 44192 15638 44220 17614
rect 44272 17128 44324 17134
rect 44272 17070 44324 17076
rect 44180 15632 44232 15638
rect 44180 15574 44232 15580
rect 44180 15156 44232 15162
rect 44180 15098 44232 15104
rect 44192 14550 44220 15098
rect 44180 14544 44232 14550
rect 44180 14486 44232 14492
rect 44180 14340 44232 14346
rect 44180 14282 44232 14288
rect 44088 12436 44140 12442
rect 44088 12378 44140 12384
rect 43996 12164 44048 12170
rect 43996 12106 44048 12112
rect 44192 12102 44220 14282
rect 44284 13530 44312 17070
rect 44362 16280 44418 16289
rect 44362 16215 44418 16224
rect 44376 15638 44404 16215
rect 44468 16046 44496 18226
rect 44548 18216 44600 18222
rect 44548 18158 44600 18164
rect 44560 17882 44588 18158
rect 44548 17876 44600 17882
rect 44548 17818 44600 17824
rect 44652 17320 44680 23054
rect 44744 22094 44772 24550
rect 44836 24070 44864 29106
rect 44928 26926 44956 30058
rect 46400 29782 46428 30194
rect 46768 29850 46796 30330
rect 47044 29850 47072 31282
rect 49252 30802 49280 56646
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 57336 54528 57388 54534
rect 57336 54470 57388 54476
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 48412 30796 48464 30802
rect 48412 30738 48464 30744
rect 49240 30796 49292 30802
rect 49240 30738 49292 30744
rect 48320 30728 48372 30734
rect 48320 30670 48372 30676
rect 48332 30326 48360 30670
rect 48320 30320 48372 30326
rect 48320 30262 48372 30268
rect 48424 29850 48452 30738
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 49516 30320 49568 30326
rect 49516 30262 49568 30268
rect 49240 30252 49292 30258
rect 49240 30194 49292 30200
rect 46756 29844 46808 29850
rect 46756 29786 46808 29792
rect 47032 29844 47084 29850
rect 47032 29786 47084 29792
rect 48412 29844 48464 29850
rect 48412 29786 48464 29792
rect 46388 29776 46440 29782
rect 46388 29718 46440 29724
rect 48136 29776 48188 29782
rect 48136 29718 48188 29724
rect 48964 29776 49016 29782
rect 48964 29718 49016 29724
rect 46112 29708 46164 29714
rect 46112 29650 46164 29656
rect 45468 29640 45520 29646
rect 45468 29582 45520 29588
rect 45192 29504 45244 29510
rect 45192 29446 45244 29452
rect 45008 28484 45060 28490
rect 45008 28426 45060 28432
rect 44916 26920 44968 26926
rect 44916 26862 44968 26868
rect 44916 26784 44968 26790
rect 44916 26726 44968 26732
rect 44928 25294 44956 26726
rect 44916 25288 44968 25294
rect 44916 25230 44968 25236
rect 44928 24886 44956 25230
rect 44916 24880 44968 24886
rect 44916 24822 44968 24828
rect 44824 24064 44876 24070
rect 44824 24006 44876 24012
rect 44744 22066 44864 22094
rect 44836 22030 44864 22066
rect 44824 22024 44876 22030
rect 44824 21966 44876 21972
rect 44836 18850 44864 21966
rect 44928 21894 44956 24822
rect 45020 23254 45048 28426
rect 45100 28076 45152 28082
rect 45100 28018 45152 28024
rect 45112 26790 45140 28018
rect 45100 26784 45152 26790
rect 45100 26726 45152 26732
rect 45204 25498 45232 29446
rect 45480 29170 45508 29582
rect 46124 29306 46152 29650
rect 46204 29640 46256 29646
rect 46204 29582 46256 29588
rect 46112 29300 46164 29306
rect 46112 29242 46164 29248
rect 45468 29164 45520 29170
rect 45468 29106 45520 29112
rect 46216 28966 46244 29582
rect 46400 29306 46428 29718
rect 47952 29572 48004 29578
rect 47952 29514 48004 29520
rect 47216 29504 47268 29510
rect 47216 29446 47268 29452
rect 46388 29300 46440 29306
rect 46388 29242 46440 29248
rect 47228 29170 47256 29446
rect 47964 29170 47992 29514
rect 47216 29164 47268 29170
rect 47216 29106 47268 29112
rect 47952 29164 48004 29170
rect 47952 29106 48004 29112
rect 46204 28960 46256 28966
rect 46204 28902 46256 28908
rect 46848 28960 46900 28966
rect 46848 28902 46900 28908
rect 46216 28762 46244 28902
rect 46204 28756 46256 28762
rect 46204 28698 46256 28704
rect 46020 28688 46072 28694
rect 46020 28630 46072 28636
rect 45652 28552 45704 28558
rect 45652 28494 45704 28500
rect 45664 28422 45692 28494
rect 45652 28416 45704 28422
rect 45652 28358 45704 28364
rect 45664 27606 45692 28358
rect 45744 28144 45796 28150
rect 45744 28086 45796 28092
rect 45652 27600 45704 27606
rect 45652 27542 45704 27548
rect 45756 27470 45784 28086
rect 45836 28076 45888 28082
rect 45836 28018 45888 28024
rect 45848 27470 45876 28018
rect 45928 27940 45980 27946
rect 45928 27882 45980 27888
rect 45940 27538 45968 27882
rect 46032 27674 46060 28630
rect 46860 28626 46888 28902
rect 47228 28762 47256 29106
rect 47216 28756 47268 28762
rect 47216 28698 47268 28704
rect 46848 28620 46900 28626
rect 46848 28562 46900 28568
rect 46664 28416 46716 28422
rect 46664 28358 46716 28364
rect 46296 28008 46348 28014
rect 46296 27950 46348 27956
rect 46020 27668 46072 27674
rect 46020 27610 46072 27616
rect 45928 27532 45980 27538
rect 45928 27474 45980 27480
rect 46308 27470 46336 27950
rect 46676 27470 46704 28358
rect 46860 28218 46888 28562
rect 46848 28212 46900 28218
rect 46848 28154 46900 28160
rect 47860 28076 47912 28082
rect 47860 28018 47912 28024
rect 47492 28008 47544 28014
rect 47492 27950 47544 27956
rect 47124 27872 47176 27878
rect 47124 27814 47176 27820
rect 45744 27464 45796 27470
rect 45744 27406 45796 27412
rect 45836 27464 45888 27470
rect 45836 27406 45888 27412
rect 46296 27464 46348 27470
rect 46296 27406 46348 27412
rect 46664 27464 46716 27470
rect 46664 27406 46716 27412
rect 45756 27130 45784 27406
rect 45744 27124 45796 27130
rect 45744 27066 45796 27072
rect 45376 26376 45428 26382
rect 45376 26318 45428 26324
rect 45388 25974 45416 26318
rect 45848 26314 45876 27406
rect 46020 26920 46072 26926
rect 46020 26862 46072 26868
rect 45928 26512 45980 26518
rect 45928 26454 45980 26460
rect 45836 26308 45888 26314
rect 45836 26250 45888 26256
rect 45376 25968 45428 25974
rect 45376 25910 45428 25916
rect 45744 25968 45796 25974
rect 45744 25910 45796 25916
rect 45192 25492 45244 25498
rect 45192 25434 45244 25440
rect 45204 24410 45232 25434
rect 45468 25152 45520 25158
rect 45468 25094 45520 25100
rect 45652 25152 45704 25158
rect 45652 25094 45704 25100
rect 45480 24818 45508 25094
rect 45468 24812 45520 24818
rect 45468 24754 45520 24760
rect 45560 24744 45612 24750
rect 45664 24698 45692 25094
rect 45612 24692 45692 24698
rect 45560 24686 45692 24692
rect 45572 24670 45692 24686
rect 45376 24608 45428 24614
rect 45376 24550 45428 24556
rect 45192 24404 45244 24410
rect 45192 24346 45244 24352
rect 45388 24138 45416 24550
rect 45376 24132 45428 24138
rect 45376 24074 45428 24080
rect 45572 23254 45600 24670
rect 45756 24614 45784 25910
rect 45836 25288 45888 25294
rect 45836 25230 45888 25236
rect 45848 24750 45876 25230
rect 45836 24744 45888 24750
rect 45836 24686 45888 24692
rect 45744 24608 45796 24614
rect 45744 24550 45796 24556
rect 45756 23322 45784 24550
rect 45744 23316 45796 23322
rect 45744 23258 45796 23264
rect 45008 23248 45060 23254
rect 45008 23190 45060 23196
rect 45560 23248 45612 23254
rect 45560 23190 45612 23196
rect 45560 23112 45612 23118
rect 45560 23054 45612 23060
rect 45572 22658 45600 23054
rect 45572 22630 45692 22658
rect 45756 22642 45784 23258
rect 45664 22574 45692 22630
rect 45744 22636 45796 22642
rect 45744 22578 45796 22584
rect 45652 22568 45704 22574
rect 45652 22510 45704 22516
rect 45560 22500 45612 22506
rect 45560 22442 45612 22448
rect 45572 22166 45600 22442
rect 45560 22160 45612 22166
rect 45560 22102 45612 22108
rect 44916 21888 44968 21894
rect 44916 21830 44968 21836
rect 45376 21888 45428 21894
rect 45376 21830 45428 21836
rect 45284 21616 45336 21622
rect 45284 21558 45336 21564
rect 45296 20806 45324 21558
rect 45284 20800 45336 20806
rect 45284 20742 45336 20748
rect 45008 19304 45060 19310
rect 45008 19246 45060 19252
rect 45020 18902 45048 19246
rect 45008 18896 45060 18902
rect 44836 18822 44956 18850
rect 45008 18838 45060 18844
rect 44824 18216 44876 18222
rect 44824 18158 44876 18164
rect 44836 17814 44864 18158
rect 44824 17808 44876 17814
rect 44824 17750 44876 17756
rect 44560 17292 44680 17320
rect 44456 16040 44508 16046
rect 44456 15982 44508 15988
rect 44364 15632 44416 15638
rect 44364 15574 44416 15580
rect 44454 15600 44510 15609
rect 44376 13938 44404 15574
rect 44454 15535 44510 15544
rect 44364 13932 44416 13938
rect 44364 13874 44416 13880
rect 44362 13696 44418 13705
rect 44362 13631 44418 13640
rect 44272 13524 44324 13530
rect 44272 13466 44324 13472
rect 44376 13462 44404 13631
rect 44364 13456 44416 13462
rect 44364 13398 44416 13404
rect 44180 12096 44232 12102
rect 44180 12038 44232 12044
rect 43996 11688 44048 11694
rect 43996 11630 44048 11636
rect 44008 11354 44036 11630
rect 43996 11348 44048 11354
rect 43996 11290 44048 11296
rect 43996 11008 44048 11014
rect 43994 10976 43996 10985
rect 44088 11008 44140 11014
rect 44048 10976 44050 10985
rect 44088 10950 44140 10956
rect 43994 10911 44050 10920
rect 44008 9994 44036 10911
rect 44100 10742 44128 10950
rect 44088 10736 44140 10742
rect 44088 10678 44140 10684
rect 44088 10464 44140 10470
rect 44088 10406 44140 10412
rect 44100 10062 44128 10406
rect 44088 10056 44140 10062
rect 44088 9998 44140 10004
rect 43996 9988 44048 9994
rect 43996 9930 44048 9936
rect 43996 9580 44048 9586
rect 43996 9522 44048 9528
rect 44008 8634 44036 9522
rect 44192 8922 44220 12038
rect 44270 11928 44326 11937
rect 44270 11863 44272 11872
rect 44324 11863 44326 11872
rect 44272 11834 44324 11840
rect 44272 10668 44324 10674
rect 44272 10610 44324 10616
rect 44284 9722 44312 10610
rect 44376 10062 44404 13398
rect 44468 11762 44496 15535
rect 44560 14958 44588 17292
rect 44640 17196 44692 17202
rect 44640 17138 44692 17144
rect 44652 15162 44680 17138
rect 44732 16584 44784 16590
rect 44732 16526 44784 16532
rect 44744 16250 44772 16526
rect 44732 16244 44784 16250
rect 44732 16186 44784 16192
rect 44928 16130 44956 18822
rect 45008 18148 45060 18154
rect 45008 18090 45060 18096
rect 44744 16102 44956 16130
rect 44640 15156 44692 15162
rect 44640 15098 44692 15104
rect 44548 14952 44600 14958
rect 44548 14894 44600 14900
rect 44548 13932 44600 13938
rect 44548 13874 44600 13880
rect 44560 13394 44588 13874
rect 44640 13728 44692 13734
rect 44640 13670 44692 13676
rect 44548 13388 44600 13394
rect 44548 13330 44600 13336
rect 44652 13326 44680 13670
rect 44640 13320 44692 13326
rect 44640 13262 44692 13268
rect 44548 12980 44600 12986
rect 44548 12922 44600 12928
rect 44560 12714 44588 12922
rect 44652 12918 44680 13262
rect 44640 12912 44692 12918
rect 44640 12854 44692 12860
rect 44548 12708 44600 12714
rect 44548 12650 44600 12656
rect 44640 12708 44692 12714
rect 44640 12650 44692 12656
rect 44456 11756 44508 11762
rect 44456 11698 44508 11704
rect 44560 11082 44588 12650
rect 44548 11076 44600 11082
rect 44548 11018 44600 11024
rect 44364 10056 44416 10062
rect 44364 9998 44416 10004
rect 44548 9988 44600 9994
rect 44548 9930 44600 9936
rect 44362 9752 44418 9761
rect 44272 9716 44324 9722
rect 44362 9687 44418 9696
rect 44272 9658 44324 9664
rect 44376 9654 44404 9687
rect 44364 9648 44416 9654
rect 44364 9590 44416 9596
rect 44192 8894 44312 8922
rect 44088 8832 44140 8838
rect 44140 8780 44220 8786
rect 44088 8774 44220 8780
rect 44100 8758 44220 8774
rect 43996 8628 44048 8634
rect 43996 8570 44048 8576
rect 44088 8492 44140 8498
rect 44088 8434 44140 8440
rect 44100 7954 44128 8434
rect 44088 7948 44140 7954
rect 44088 7890 44140 7896
rect 44088 7744 44140 7750
rect 44088 7686 44140 7692
rect 43996 7472 44048 7478
rect 43996 7414 44048 7420
rect 43902 6896 43958 6905
rect 43902 6831 43958 6840
rect 43916 6730 43944 6831
rect 43904 6724 43956 6730
rect 43904 6666 43956 6672
rect 43916 6458 43944 6666
rect 43904 6452 43956 6458
rect 43904 6394 43956 6400
rect 44008 5574 44036 7414
rect 44100 7410 44128 7686
rect 44192 7410 44220 8758
rect 44284 7886 44312 8894
rect 44560 8430 44588 9930
rect 44652 8838 44680 12650
rect 44744 9586 44772 16102
rect 44824 15632 44876 15638
rect 44824 15574 44876 15580
rect 44836 15026 44864 15574
rect 44914 15056 44970 15065
rect 44824 15020 44876 15026
rect 44914 14991 44916 15000
rect 44824 14962 44876 14968
rect 44968 14991 44970 15000
rect 44916 14962 44968 14968
rect 44836 13870 44864 14962
rect 44928 14618 44956 14962
rect 44916 14612 44968 14618
rect 44916 14554 44968 14560
rect 44824 13864 44876 13870
rect 44824 13806 44876 13812
rect 44928 12986 44956 14554
rect 45020 13569 45048 18090
rect 45284 17672 45336 17678
rect 45284 17614 45336 17620
rect 45100 17604 45152 17610
rect 45100 17546 45152 17552
rect 45112 16998 45140 17546
rect 45296 17105 45324 17614
rect 45282 17096 45338 17105
rect 45282 17031 45338 17040
rect 45100 16992 45152 16998
rect 45100 16934 45152 16940
rect 45006 13560 45062 13569
rect 45006 13495 45062 13504
rect 44916 12980 44968 12986
rect 44916 12922 44968 12928
rect 44928 12714 44956 12922
rect 44916 12708 44968 12714
rect 44916 12650 44968 12656
rect 44916 12368 44968 12374
rect 44916 12310 44968 12316
rect 44928 11762 44956 12310
rect 45020 12209 45048 13495
rect 45006 12200 45062 12209
rect 45006 12135 45062 12144
rect 44916 11756 44968 11762
rect 44916 11698 44968 11704
rect 45112 11626 45140 16934
rect 45388 16522 45416 21830
rect 45572 20890 45600 22102
rect 45664 22094 45692 22510
rect 45664 22066 45784 22094
rect 45756 22030 45784 22066
rect 45744 22024 45796 22030
rect 45744 21966 45796 21972
rect 45756 21146 45784 21966
rect 45744 21140 45796 21146
rect 45744 21082 45796 21088
rect 45572 20862 45784 20890
rect 45756 20806 45784 20862
rect 45744 20800 45796 20806
rect 45744 20742 45796 20748
rect 45560 20460 45612 20466
rect 45560 20402 45612 20408
rect 45572 19854 45600 20402
rect 45756 20398 45784 20742
rect 45744 20392 45796 20398
rect 45744 20334 45796 20340
rect 45756 19854 45784 20334
rect 45560 19848 45612 19854
rect 45560 19790 45612 19796
rect 45744 19848 45796 19854
rect 45744 19790 45796 19796
rect 45652 19780 45704 19786
rect 45652 19722 45704 19728
rect 45664 18290 45692 19722
rect 45756 19446 45784 19790
rect 45744 19440 45796 19446
rect 45744 19382 45796 19388
rect 45756 18834 45784 19382
rect 45848 19174 45876 24686
rect 45940 22094 45968 26454
rect 46032 26382 46060 26862
rect 46112 26784 46164 26790
rect 46112 26726 46164 26732
rect 46124 26586 46152 26726
rect 46112 26580 46164 26586
rect 46112 26522 46164 26528
rect 46204 26512 46256 26518
rect 46204 26454 46256 26460
rect 46020 26376 46072 26382
rect 46020 26318 46072 26324
rect 46032 25702 46060 26318
rect 46112 25832 46164 25838
rect 46112 25774 46164 25780
rect 46020 25696 46072 25702
rect 46020 25638 46072 25644
rect 46032 25498 46060 25638
rect 46020 25492 46072 25498
rect 46020 25434 46072 25440
rect 46032 24750 46060 25434
rect 46020 24744 46072 24750
rect 46020 24686 46072 24692
rect 46032 23866 46060 24686
rect 46020 23860 46072 23866
rect 46020 23802 46072 23808
rect 46032 23118 46060 23802
rect 46020 23112 46072 23118
rect 46020 23054 46072 23060
rect 46032 22778 46060 23054
rect 46020 22772 46072 22778
rect 46020 22714 46072 22720
rect 46124 22574 46152 25774
rect 46216 25362 46244 26454
rect 46204 25356 46256 25362
rect 46204 25298 46256 25304
rect 46216 24818 46244 25298
rect 46204 24812 46256 24818
rect 46204 24754 46256 24760
rect 46216 23798 46244 24754
rect 46204 23792 46256 23798
rect 46204 23734 46256 23740
rect 46204 22636 46256 22642
rect 46204 22578 46256 22584
rect 46112 22568 46164 22574
rect 46110 22536 46112 22545
rect 46164 22536 46166 22545
rect 46110 22471 46166 22480
rect 45940 22066 46060 22094
rect 46032 19922 46060 22066
rect 46020 19916 46072 19922
rect 46020 19858 46072 19864
rect 46020 19372 46072 19378
rect 46020 19314 46072 19320
rect 45836 19168 45888 19174
rect 45836 19110 45888 19116
rect 46032 18970 46060 19314
rect 46020 18964 46072 18970
rect 46020 18906 46072 18912
rect 45744 18828 45796 18834
rect 45744 18770 45796 18776
rect 45756 18630 45784 18770
rect 45744 18624 45796 18630
rect 45744 18566 45796 18572
rect 45928 18624 45980 18630
rect 45928 18566 45980 18572
rect 45652 18284 45704 18290
rect 45652 18226 45704 18232
rect 45756 17785 45784 18566
rect 45742 17776 45798 17785
rect 45742 17711 45798 17720
rect 45468 17672 45520 17678
rect 45466 17640 45468 17649
rect 45744 17672 45796 17678
rect 45520 17640 45522 17649
rect 45744 17614 45796 17620
rect 45466 17575 45522 17584
rect 45652 17264 45704 17270
rect 45652 17206 45704 17212
rect 45560 17060 45612 17066
rect 45560 17002 45612 17008
rect 45468 16992 45520 16998
rect 45468 16934 45520 16940
rect 45480 16794 45508 16934
rect 45468 16788 45520 16794
rect 45468 16730 45520 16736
rect 45376 16516 45428 16522
rect 45376 16458 45428 16464
rect 45192 16176 45244 16182
rect 45192 16118 45244 16124
rect 45204 15881 45232 16118
rect 45572 16114 45600 17002
rect 45560 16108 45612 16114
rect 45560 16050 45612 16056
rect 45190 15872 45246 15881
rect 45664 15858 45692 17206
rect 45756 16114 45784 17614
rect 45940 17202 45968 18566
rect 46020 17876 46072 17882
rect 46020 17818 46072 17824
rect 46032 17610 46060 17818
rect 46112 17808 46164 17814
rect 46112 17750 46164 17756
rect 46020 17604 46072 17610
rect 46020 17546 46072 17552
rect 46124 17338 46152 17750
rect 46112 17332 46164 17338
rect 46032 17292 46112 17320
rect 45928 17196 45980 17202
rect 45928 17138 45980 17144
rect 45926 16144 45982 16153
rect 45744 16108 45796 16114
rect 46032 16114 46060 17292
rect 46112 17274 46164 17280
rect 46112 17060 46164 17066
rect 46112 17002 46164 17008
rect 46124 16590 46152 17002
rect 46112 16584 46164 16590
rect 46112 16526 46164 16532
rect 46124 16425 46152 16526
rect 46110 16416 46166 16425
rect 46110 16351 46166 16360
rect 46216 16250 46244 22578
rect 46308 22166 46336 27406
rect 46572 26988 46624 26994
rect 46572 26930 46624 26936
rect 46584 26450 46612 26930
rect 46676 26790 46704 27406
rect 47136 27062 47164 27814
rect 47216 27668 47268 27674
rect 47216 27610 47268 27616
rect 47124 27056 47176 27062
rect 47124 26998 47176 27004
rect 46664 26784 46716 26790
rect 46664 26726 46716 26732
rect 47032 26580 47084 26586
rect 47032 26522 47084 26528
rect 46572 26444 46624 26450
rect 46572 26386 46624 26392
rect 46584 25906 46612 26386
rect 46940 26376 46992 26382
rect 46940 26318 46992 26324
rect 46952 25906 46980 26318
rect 46572 25900 46624 25906
rect 46572 25842 46624 25848
rect 46940 25900 46992 25906
rect 46940 25842 46992 25848
rect 46584 24818 46612 25842
rect 47044 25838 47072 26522
rect 47136 26314 47164 26998
rect 47228 26586 47256 27610
rect 47504 27538 47532 27950
rect 47872 27606 47900 28018
rect 47964 27606 47992 29106
rect 48148 28966 48176 29718
rect 48976 29102 49004 29718
rect 49252 29714 49280 30194
rect 49424 30048 49476 30054
rect 49424 29990 49476 29996
rect 49240 29708 49292 29714
rect 49240 29650 49292 29656
rect 49252 29170 49280 29650
rect 49240 29164 49292 29170
rect 49240 29106 49292 29112
rect 48964 29096 49016 29102
rect 48964 29038 49016 29044
rect 49332 29096 49384 29102
rect 49332 29038 49384 29044
rect 48136 28960 48188 28966
rect 48136 28902 48188 28908
rect 49344 28626 49372 29038
rect 49332 28620 49384 28626
rect 49332 28562 49384 28568
rect 49436 28558 49464 29990
rect 49528 29170 49556 30262
rect 50988 29640 51040 29646
rect 50908 29588 50988 29594
rect 50908 29582 51040 29588
rect 51816 29640 51868 29646
rect 51816 29582 51868 29588
rect 50908 29566 51028 29582
rect 50908 29458 50936 29566
rect 50816 29430 50936 29458
rect 50988 29504 51040 29510
rect 50988 29446 51040 29452
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 49608 29300 49660 29306
rect 49608 29242 49660 29248
rect 49516 29164 49568 29170
rect 49516 29106 49568 29112
rect 49620 28558 49648 29242
rect 49792 29164 49844 29170
rect 49792 29106 49844 29112
rect 49424 28552 49476 28558
rect 49424 28494 49476 28500
rect 49608 28552 49660 28558
rect 49608 28494 49660 28500
rect 48504 28076 48556 28082
rect 48504 28018 48556 28024
rect 47860 27600 47912 27606
rect 47860 27542 47912 27548
rect 47952 27600 48004 27606
rect 47952 27542 48004 27548
rect 47492 27532 47544 27538
rect 47492 27474 47544 27480
rect 47308 27464 47360 27470
rect 47308 27406 47360 27412
rect 47320 27130 47348 27406
rect 47308 27124 47360 27130
rect 47308 27066 47360 27072
rect 47216 26580 47268 26586
rect 47216 26522 47268 26528
rect 47124 26308 47176 26314
rect 47124 26250 47176 26256
rect 47032 25832 47084 25838
rect 47032 25774 47084 25780
rect 47136 25770 47164 26250
rect 47124 25764 47176 25770
rect 47124 25706 47176 25712
rect 47504 25498 47532 27474
rect 48516 27130 48544 28018
rect 49424 28008 49476 28014
rect 49424 27950 49476 27956
rect 49436 27470 49464 27950
rect 49620 27674 49648 28494
rect 49804 28490 49832 29106
rect 50816 28694 50844 29430
rect 50896 29232 50948 29238
rect 50896 29174 50948 29180
rect 50804 28688 50856 28694
rect 50804 28630 50856 28636
rect 49792 28484 49844 28490
rect 49792 28426 49844 28432
rect 49700 28076 49752 28082
rect 49700 28018 49752 28024
rect 49608 27668 49660 27674
rect 49608 27610 49660 27616
rect 49712 27470 49740 28018
rect 49804 28014 49832 28426
rect 50068 28416 50120 28422
rect 50068 28358 50120 28364
rect 49792 28008 49844 28014
rect 49792 27950 49844 27956
rect 50080 27713 50108 28358
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50816 28082 50844 28630
rect 50620 28076 50672 28082
rect 50620 28018 50672 28024
rect 50804 28076 50856 28082
rect 50804 28018 50856 28024
rect 50066 27704 50122 27713
rect 50066 27639 50122 27648
rect 50632 27470 50660 28018
rect 50908 27826 50936 29174
rect 51000 28966 51028 29446
rect 51828 29306 51856 29582
rect 51816 29300 51868 29306
rect 51816 29242 51868 29248
rect 51172 29164 51224 29170
rect 51172 29106 51224 29112
rect 54116 29164 54168 29170
rect 54116 29106 54168 29112
rect 55220 29164 55272 29170
rect 55220 29106 55272 29112
rect 50988 28960 51040 28966
rect 50988 28902 51040 28908
rect 51000 28626 51028 28902
rect 50988 28620 51040 28626
rect 50988 28562 51040 28568
rect 51000 27946 51028 28562
rect 51184 28490 51212 29106
rect 53932 28620 53984 28626
rect 53932 28562 53984 28568
rect 51356 28552 51408 28558
rect 51356 28494 51408 28500
rect 52920 28552 52972 28558
rect 52920 28494 52972 28500
rect 53748 28552 53800 28558
rect 53748 28494 53800 28500
rect 51172 28484 51224 28490
rect 51172 28426 51224 28432
rect 51080 28008 51132 28014
rect 51184 27996 51212 28426
rect 51368 28082 51396 28494
rect 51356 28076 51408 28082
rect 51356 28018 51408 28024
rect 52828 28076 52880 28082
rect 52932 28064 52960 28494
rect 53012 28416 53064 28422
rect 53012 28358 53064 28364
rect 53024 28082 53052 28358
rect 53760 28082 53788 28494
rect 53840 28416 53892 28422
rect 53840 28358 53892 28364
rect 52880 28036 52960 28064
rect 52828 28018 52880 28024
rect 51132 27968 51212 27996
rect 51080 27950 51132 27956
rect 50988 27940 51040 27946
rect 50988 27882 51040 27888
rect 50908 27798 51028 27826
rect 49424 27464 49476 27470
rect 49424 27406 49476 27412
rect 49700 27464 49752 27470
rect 49700 27406 49752 27412
rect 50620 27464 50672 27470
rect 50620 27406 50672 27412
rect 50896 27464 50948 27470
rect 50896 27406 50948 27412
rect 49516 27328 49568 27334
rect 49516 27270 49568 27276
rect 48504 27124 48556 27130
rect 48504 27066 48556 27072
rect 47584 27056 47636 27062
rect 47584 26998 47636 27004
rect 47596 26382 47624 26998
rect 48044 26988 48096 26994
rect 48044 26930 48096 26936
rect 48136 26988 48188 26994
rect 48136 26930 48188 26936
rect 49240 26988 49292 26994
rect 49240 26930 49292 26936
rect 47952 26920 48004 26926
rect 47952 26862 48004 26868
rect 47964 26450 47992 26862
rect 48056 26518 48084 26930
rect 48044 26512 48096 26518
rect 48044 26454 48096 26460
rect 47952 26444 48004 26450
rect 47952 26386 48004 26392
rect 47584 26376 47636 26382
rect 48148 26330 48176 26930
rect 48228 26852 48280 26858
rect 48228 26794 48280 26800
rect 48240 26518 48268 26794
rect 48780 26784 48832 26790
rect 48780 26726 48832 26732
rect 48228 26512 48280 26518
rect 48228 26454 48280 26460
rect 48792 26382 48820 26726
rect 49252 26382 49280 26930
rect 49528 26382 49556 27270
rect 49712 26586 49740 27406
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50632 26790 50660 27406
rect 50712 27328 50764 27334
rect 50712 27270 50764 27276
rect 50724 27062 50752 27270
rect 50908 27062 50936 27406
rect 50712 27056 50764 27062
rect 50896 27056 50948 27062
rect 50712 26998 50764 27004
rect 50816 27004 50896 27010
rect 50816 26998 50948 27004
rect 50620 26784 50672 26790
rect 50620 26726 50672 26732
rect 49700 26580 49752 26586
rect 49700 26522 49752 26528
rect 50632 26382 50660 26726
rect 50724 26382 50752 26998
rect 50816 26982 50936 26998
rect 47584 26318 47636 26324
rect 47492 25492 47544 25498
rect 47492 25434 47544 25440
rect 47308 25356 47360 25362
rect 47308 25298 47360 25304
rect 47124 25220 47176 25226
rect 47124 25162 47176 25168
rect 47136 24886 47164 25162
rect 47320 24954 47348 25298
rect 47308 24948 47360 24954
rect 47308 24890 47360 24896
rect 47124 24880 47176 24886
rect 47124 24822 47176 24828
rect 46572 24812 46624 24818
rect 46572 24754 46624 24760
rect 46584 22642 46612 24754
rect 47136 24410 47164 24822
rect 47124 24404 47176 24410
rect 47124 24346 47176 24352
rect 46664 24200 46716 24206
rect 46848 24200 46900 24206
rect 46664 24142 46716 24148
rect 46768 24148 46848 24154
rect 46768 24142 46900 24148
rect 46676 23730 46704 24142
rect 46768 24126 46888 24142
rect 46940 24132 46992 24138
rect 46768 23730 46796 24126
rect 46940 24074 46992 24080
rect 46848 24064 46900 24070
rect 46848 24006 46900 24012
rect 46860 23866 46888 24006
rect 46848 23860 46900 23866
rect 46848 23802 46900 23808
rect 46952 23730 46980 24074
rect 46664 23724 46716 23730
rect 46664 23666 46716 23672
rect 46756 23724 46808 23730
rect 46756 23666 46808 23672
rect 46940 23724 46992 23730
rect 46940 23666 46992 23672
rect 47308 23724 47360 23730
rect 47308 23666 47360 23672
rect 46676 23322 46704 23666
rect 46664 23316 46716 23322
rect 46664 23258 46716 23264
rect 46768 23118 46796 23666
rect 46756 23112 46808 23118
rect 46756 23054 46808 23060
rect 46664 22772 46716 22778
rect 46664 22714 46716 22720
rect 46572 22636 46624 22642
rect 46572 22578 46624 22584
rect 46296 22160 46348 22166
rect 46296 22102 46348 22108
rect 46584 21894 46612 22578
rect 46572 21888 46624 21894
rect 46572 21830 46624 21836
rect 46584 21622 46612 21830
rect 46572 21616 46624 21622
rect 46572 21558 46624 21564
rect 46296 19984 46348 19990
rect 46296 19926 46348 19932
rect 46308 19310 46336 19926
rect 46296 19304 46348 19310
rect 46296 19246 46348 19252
rect 46204 16244 46256 16250
rect 46204 16186 46256 16192
rect 45926 16079 45982 16088
rect 46020 16108 46072 16114
rect 45744 16050 45796 16056
rect 45836 16040 45888 16046
rect 45836 15982 45888 15988
rect 45190 15807 45246 15816
rect 45572 15830 45692 15858
rect 45376 15564 45428 15570
rect 45376 15506 45428 15512
rect 45388 15473 45416 15506
rect 45374 15464 45430 15473
rect 45374 15399 45430 15408
rect 45284 15360 45336 15366
rect 45282 15328 45284 15337
rect 45336 15328 45338 15337
rect 45572 15314 45600 15830
rect 45848 15706 45876 15982
rect 45744 15700 45796 15706
rect 45744 15642 45796 15648
rect 45836 15700 45888 15706
rect 45836 15642 45888 15648
rect 45756 15366 45784 15642
rect 45282 15263 45338 15272
rect 45388 15286 45600 15314
rect 45652 15360 45704 15366
rect 45652 15302 45704 15308
rect 45744 15360 45796 15366
rect 45796 15320 45876 15348
rect 45744 15302 45796 15308
rect 45192 15156 45244 15162
rect 45192 15098 45244 15104
rect 45204 15026 45232 15098
rect 45192 15020 45244 15026
rect 45192 14962 45244 14968
rect 45282 14920 45338 14929
rect 45282 14855 45338 14864
rect 45296 14056 45324 14855
rect 45388 14346 45416 15286
rect 45664 15026 45692 15302
rect 45652 15020 45704 15026
rect 45652 14962 45704 14968
rect 45744 15020 45796 15026
rect 45744 14962 45796 14968
rect 45468 14884 45520 14890
rect 45468 14826 45520 14832
rect 45560 14884 45612 14890
rect 45560 14826 45612 14832
rect 45376 14340 45428 14346
rect 45376 14282 45428 14288
rect 45204 14028 45416 14056
rect 45204 13190 45232 14028
rect 45388 13938 45416 14028
rect 45284 13932 45336 13938
rect 45284 13874 45336 13880
rect 45376 13932 45428 13938
rect 45376 13874 45428 13880
rect 45192 13184 45244 13190
rect 45192 13126 45244 13132
rect 45192 12776 45244 12782
rect 45192 12718 45244 12724
rect 45204 11937 45232 12718
rect 45296 12374 45324 13874
rect 45376 13320 45428 13326
rect 45376 13262 45428 13268
rect 45388 13161 45416 13262
rect 45374 13152 45430 13161
rect 45374 13087 45430 13096
rect 45376 12844 45428 12850
rect 45376 12786 45428 12792
rect 45284 12368 45336 12374
rect 45284 12310 45336 12316
rect 45284 12164 45336 12170
rect 45284 12106 45336 12112
rect 45190 11928 45246 11937
rect 45190 11863 45246 11872
rect 45100 11620 45152 11626
rect 45100 11562 45152 11568
rect 45100 11280 45152 11286
rect 45100 11222 45152 11228
rect 44824 11144 44876 11150
rect 44824 11086 44876 11092
rect 44732 9580 44784 9586
rect 44732 9522 44784 9528
rect 44836 9353 44864 11086
rect 44822 9344 44878 9353
rect 44822 9279 44878 9288
rect 44836 8974 44864 9279
rect 45112 9110 45140 11222
rect 45296 10033 45324 12106
rect 45388 12084 45416 12786
rect 45480 12322 45508 14826
rect 45572 14618 45600 14826
rect 45560 14612 45612 14618
rect 45560 14554 45612 14560
rect 45652 14612 45704 14618
rect 45756 14600 45784 14962
rect 45704 14572 45784 14600
rect 45652 14554 45704 14560
rect 45848 14550 45876 15320
rect 45940 15162 45968 16079
rect 46020 16050 46072 16056
rect 46204 16108 46256 16114
rect 46204 16050 46256 16056
rect 46112 15904 46164 15910
rect 46112 15846 46164 15852
rect 46124 15570 46152 15846
rect 46112 15564 46164 15570
rect 46112 15506 46164 15512
rect 46216 15473 46244 16050
rect 46202 15464 46258 15473
rect 46202 15399 46258 15408
rect 46204 15360 46256 15366
rect 46204 15302 46256 15308
rect 45928 15156 45980 15162
rect 45928 15098 45980 15104
rect 45940 15026 45968 15098
rect 46216 15094 46244 15302
rect 46204 15088 46256 15094
rect 46204 15030 46256 15036
rect 45928 15020 45980 15026
rect 46112 15020 46164 15026
rect 45928 14962 45980 14968
rect 46032 14980 46112 15008
rect 45928 14816 45980 14822
rect 45928 14758 45980 14764
rect 45836 14544 45888 14550
rect 45836 14486 45888 14492
rect 45652 14408 45704 14414
rect 45558 14376 45614 14385
rect 45652 14350 45704 14356
rect 45558 14311 45614 14320
rect 45572 14278 45600 14311
rect 45560 14272 45612 14278
rect 45560 14214 45612 14220
rect 45664 13258 45692 14350
rect 45744 14272 45796 14278
rect 45744 14214 45796 14220
rect 45756 13433 45784 14214
rect 45940 14074 45968 14758
rect 46032 14618 46060 14980
rect 46112 14962 46164 14968
rect 46308 14906 46336 19246
rect 46388 18828 46440 18834
rect 46388 18770 46440 18776
rect 46400 18358 46428 18770
rect 46388 18352 46440 18358
rect 46388 18294 46440 18300
rect 46388 17672 46440 17678
rect 46388 17614 46440 17620
rect 46480 17650 46532 17656
rect 46400 17338 46428 17614
rect 46480 17592 46532 17598
rect 46388 17332 46440 17338
rect 46388 17274 46440 17280
rect 46492 16674 46520 17592
rect 46676 17218 46704 22714
rect 46768 22710 46796 23054
rect 47320 22710 47348 23666
rect 46756 22704 46808 22710
rect 46756 22646 46808 22652
rect 47308 22704 47360 22710
rect 47308 22646 47360 22652
rect 47124 22024 47176 22030
rect 47124 21966 47176 21972
rect 46940 21344 46992 21350
rect 46938 21312 46940 21321
rect 46992 21312 46994 21321
rect 46938 21247 46994 21256
rect 46952 21146 46980 21247
rect 46940 21140 46992 21146
rect 46940 21082 46992 21088
rect 47136 20058 47164 21966
rect 47124 20052 47176 20058
rect 47124 19994 47176 20000
rect 46756 19304 46808 19310
rect 46756 19246 46808 19252
rect 46768 18766 46796 19246
rect 46756 18760 46808 18766
rect 46756 18702 46808 18708
rect 46940 18760 46992 18766
rect 46940 18702 46992 18708
rect 46848 17536 46900 17542
rect 46848 17478 46900 17484
rect 46860 17338 46888 17478
rect 46848 17332 46900 17338
rect 46848 17274 46900 17280
rect 46124 14878 46336 14906
rect 46400 16646 46520 16674
rect 46584 17190 46704 17218
rect 46020 14612 46072 14618
rect 46020 14554 46072 14560
rect 45928 14068 45980 14074
rect 45928 14010 45980 14016
rect 45836 13932 45888 13938
rect 45836 13874 45888 13880
rect 45742 13424 45798 13433
rect 45742 13359 45798 13368
rect 45652 13252 45704 13258
rect 45652 13194 45704 13200
rect 45480 12306 45600 12322
rect 45480 12300 45612 12306
rect 45480 12294 45560 12300
rect 45560 12242 45612 12248
rect 45468 12232 45520 12238
rect 45466 12200 45468 12209
rect 45520 12200 45522 12209
rect 45664 12170 45692 13194
rect 45466 12135 45522 12144
rect 45652 12164 45704 12170
rect 45652 12106 45704 12112
rect 45468 12096 45520 12102
rect 45388 12056 45468 12084
rect 45468 12038 45520 12044
rect 45560 12096 45612 12102
rect 45560 12038 45612 12044
rect 45376 10464 45428 10470
rect 45376 10406 45428 10412
rect 45388 10198 45416 10406
rect 45376 10192 45428 10198
rect 45376 10134 45428 10140
rect 45282 10024 45338 10033
rect 45282 9959 45338 9968
rect 45296 9586 45324 9959
rect 45480 9722 45508 12038
rect 45572 11898 45600 12038
rect 45650 11928 45706 11937
rect 45560 11892 45612 11898
rect 45650 11863 45706 11872
rect 45560 11834 45612 11840
rect 45560 11756 45612 11762
rect 45560 11698 45612 11704
rect 45572 11218 45600 11698
rect 45664 11626 45692 11863
rect 45652 11620 45704 11626
rect 45652 11562 45704 11568
rect 45560 11212 45612 11218
rect 45560 11154 45612 11160
rect 45558 11112 45614 11121
rect 45558 11047 45614 11056
rect 45572 10742 45600 11047
rect 45560 10736 45612 10742
rect 45560 10678 45612 10684
rect 45468 9716 45520 9722
rect 45468 9658 45520 9664
rect 45284 9580 45336 9586
rect 45284 9522 45336 9528
rect 45100 9104 45152 9110
rect 45100 9046 45152 9052
rect 44916 9036 44968 9042
rect 44916 8978 44968 8984
rect 44824 8968 44876 8974
rect 44824 8910 44876 8916
rect 44640 8832 44692 8838
rect 44640 8774 44692 8780
rect 44928 8498 44956 8978
rect 45296 8974 45324 9522
rect 45572 9518 45600 10678
rect 45664 10606 45692 11562
rect 45756 11540 45784 13359
rect 45848 12753 45876 13874
rect 46032 13462 46060 14554
rect 45928 13456 45980 13462
rect 45928 13398 45980 13404
rect 46020 13456 46072 13462
rect 46020 13398 46072 13404
rect 45940 12986 45968 13398
rect 45928 12980 45980 12986
rect 45928 12922 45980 12928
rect 46032 12918 46060 13398
rect 46020 12912 46072 12918
rect 46020 12854 46072 12860
rect 45834 12744 45890 12753
rect 45834 12679 45890 12688
rect 46124 12442 46152 14878
rect 46296 14544 46348 14550
rect 46296 14486 46348 14492
rect 46308 14362 46336 14486
rect 46216 14334 46336 14362
rect 46216 13938 46244 14334
rect 46296 14272 46348 14278
rect 46296 14214 46348 14220
rect 46204 13932 46256 13938
rect 46204 13874 46256 13880
rect 46202 13288 46258 13297
rect 46202 13223 46258 13232
rect 46216 13190 46244 13223
rect 46204 13184 46256 13190
rect 46204 13126 46256 13132
rect 46202 12744 46258 12753
rect 46202 12679 46258 12688
rect 46112 12436 46164 12442
rect 46112 12378 46164 12384
rect 45928 12300 45980 12306
rect 45928 12242 45980 12248
rect 45940 11898 45968 12242
rect 46112 12164 46164 12170
rect 46112 12106 46164 12112
rect 45928 11892 45980 11898
rect 45928 11834 45980 11840
rect 46124 11762 46152 12106
rect 46216 11762 46244 12679
rect 46308 12170 46336 14214
rect 46400 13530 46428 16646
rect 46480 16584 46532 16590
rect 46480 16526 46532 16532
rect 46388 13524 46440 13530
rect 46388 13466 46440 13472
rect 46388 13388 46440 13394
rect 46388 13330 46440 13336
rect 46400 12646 46428 13330
rect 46388 12640 46440 12646
rect 46388 12582 46440 12588
rect 46386 12200 46442 12209
rect 46296 12164 46348 12170
rect 46386 12135 46442 12144
rect 46296 12106 46348 12112
rect 46296 11892 46348 11898
rect 46296 11834 46348 11840
rect 46112 11756 46164 11762
rect 46112 11698 46164 11704
rect 46204 11756 46256 11762
rect 46204 11698 46256 11704
rect 45756 11512 46060 11540
rect 45928 11280 45980 11286
rect 45928 11222 45980 11228
rect 45744 11076 45796 11082
rect 45796 11036 45876 11064
rect 45744 11018 45796 11024
rect 45742 10840 45798 10849
rect 45742 10775 45798 10784
rect 45652 10600 45704 10606
rect 45652 10542 45704 10548
rect 45652 10260 45704 10266
rect 45652 10202 45704 10208
rect 45560 9512 45612 9518
rect 45560 9454 45612 9460
rect 45284 8968 45336 8974
rect 45284 8910 45336 8916
rect 44916 8492 44968 8498
rect 44916 8434 44968 8440
rect 44456 8424 44508 8430
rect 44456 8366 44508 8372
rect 44548 8424 44600 8430
rect 44548 8366 44600 8372
rect 44468 7886 44496 8366
rect 44272 7880 44324 7886
rect 44272 7822 44324 7828
rect 44456 7880 44508 7886
rect 44560 7857 44588 8366
rect 44456 7822 44508 7828
rect 44546 7848 44602 7857
rect 44468 7546 44496 7822
rect 44546 7783 44548 7792
rect 44600 7783 44602 7792
rect 44548 7754 44600 7760
rect 44560 7723 44588 7754
rect 44456 7540 44508 7546
rect 44456 7482 44508 7488
rect 44928 7410 44956 8434
rect 45296 8378 45324 8910
rect 45572 8906 45600 9454
rect 45664 8945 45692 10202
rect 45756 10062 45784 10775
rect 45848 10470 45876 11036
rect 45940 11014 45968 11222
rect 45928 11008 45980 11014
rect 45928 10950 45980 10956
rect 45836 10464 45888 10470
rect 45836 10406 45888 10412
rect 45926 10296 45982 10305
rect 45926 10231 45928 10240
rect 45980 10231 45982 10240
rect 45928 10202 45980 10208
rect 45744 10056 45796 10062
rect 45744 9998 45796 10004
rect 45928 9988 45980 9994
rect 45928 9930 45980 9936
rect 45744 9920 45796 9926
rect 45744 9862 45796 9868
rect 45650 8936 45706 8945
rect 45560 8900 45612 8906
rect 45650 8871 45706 8880
rect 45560 8842 45612 8848
rect 45374 8528 45430 8537
rect 45374 8463 45376 8472
rect 45428 8463 45430 8472
rect 45376 8434 45428 8440
rect 45572 8430 45600 8842
rect 45650 8800 45706 8809
rect 45650 8735 45706 8744
rect 45204 8350 45324 8378
rect 45560 8424 45612 8430
rect 45560 8366 45612 8372
rect 44088 7404 44140 7410
rect 44088 7346 44140 7352
rect 44180 7404 44232 7410
rect 44180 7346 44232 7352
rect 44916 7404 44968 7410
rect 44916 7346 44968 7352
rect 44272 7268 44324 7274
rect 44272 7210 44324 7216
rect 44284 5642 44312 7210
rect 44364 7200 44416 7206
rect 44364 7142 44416 7148
rect 44376 6730 44404 7142
rect 44364 6724 44416 6730
rect 44364 6666 44416 6672
rect 44928 6254 44956 7346
rect 45008 6452 45060 6458
rect 45008 6394 45060 6400
rect 44916 6248 44968 6254
rect 44916 6190 44968 6196
rect 44640 6112 44692 6118
rect 44640 6054 44692 6060
rect 44272 5636 44324 5642
rect 44272 5578 44324 5584
rect 43996 5568 44048 5574
rect 43996 5510 44048 5516
rect 44652 5234 44680 6054
rect 44928 5642 44956 6190
rect 44916 5636 44968 5642
rect 44916 5578 44968 5584
rect 44640 5228 44692 5234
rect 44640 5170 44692 5176
rect 44454 4720 44510 4729
rect 44454 4655 44510 4664
rect 44180 4480 44232 4486
rect 44180 4422 44232 4428
rect 43812 3528 43864 3534
rect 43812 3470 43864 3476
rect 43720 3460 43772 3466
rect 43720 3402 43772 3408
rect 43732 3194 43760 3402
rect 44192 3398 44220 4422
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 43720 3188 43772 3194
rect 43720 3130 43772 3136
rect 43536 2576 43588 2582
rect 43536 2518 43588 2524
rect 42248 2508 42300 2514
rect 42248 2450 42300 2456
rect 43548 2378 43576 2518
rect 40684 2372 40736 2378
rect 40684 2314 40736 2320
rect 43536 2372 43588 2378
rect 43536 2314 43588 2320
rect 38660 2304 38712 2310
rect 38660 2246 38712 2252
rect 38568 2032 38620 2038
rect 38568 1974 38620 1980
rect 38672 800 38700 2246
rect 44468 800 44496 4655
rect 45020 4214 45048 6394
rect 45204 4865 45232 8350
rect 45284 8288 45336 8294
rect 45284 8230 45336 8236
rect 45296 7206 45324 8230
rect 45284 7200 45336 7206
rect 45284 7142 45336 7148
rect 45560 6996 45612 7002
rect 45560 6938 45612 6944
rect 45376 6860 45428 6866
rect 45376 6802 45428 6808
rect 45284 6724 45336 6730
rect 45284 6666 45336 6672
rect 45296 5778 45324 6666
rect 45284 5772 45336 5778
rect 45284 5714 45336 5720
rect 45284 5228 45336 5234
rect 45284 5170 45336 5176
rect 45190 4856 45246 4865
rect 45190 4791 45246 4800
rect 45204 4690 45232 4791
rect 45192 4684 45244 4690
rect 45192 4626 45244 4632
rect 45192 4548 45244 4554
rect 45192 4490 45244 4496
rect 45008 4208 45060 4214
rect 45008 4150 45060 4156
rect 45204 2650 45232 4490
rect 45296 4146 45324 5170
rect 45284 4140 45336 4146
rect 45284 4082 45336 4088
rect 45296 3602 45324 4082
rect 45284 3596 45336 3602
rect 45284 3538 45336 3544
rect 45296 3126 45324 3538
rect 45388 3126 45416 6802
rect 45468 5704 45520 5710
rect 45468 5646 45520 5652
rect 45480 5114 45508 5646
rect 45572 5302 45600 6938
rect 45664 5642 45692 8735
rect 45756 7546 45784 9862
rect 45940 9654 45968 9930
rect 45928 9648 45980 9654
rect 45834 9616 45890 9625
rect 45928 9590 45980 9596
rect 45834 9551 45836 9560
rect 45888 9551 45890 9560
rect 45836 9522 45888 9528
rect 45940 9042 45968 9590
rect 46032 9586 46060 11512
rect 46124 11121 46152 11698
rect 46308 11642 46336 11834
rect 46216 11614 46336 11642
rect 46110 11112 46166 11121
rect 46110 11047 46166 11056
rect 46112 10668 46164 10674
rect 46112 10610 46164 10616
rect 46124 10266 46152 10610
rect 46112 10260 46164 10266
rect 46112 10202 46164 10208
rect 46216 9994 46244 11614
rect 46296 10668 46348 10674
rect 46296 10610 46348 10616
rect 46204 9988 46256 9994
rect 46204 9930 46256 9936
rect 46020 9580 46072 9586
rect 46020 9522 46072 9528
rect 46032 9042 46060 9522
rect 46204 9512 46256 9518
rect 46308 9489 46336 10610
rect 46204 9454 46256 9460
rect 46294 9480 46350 9489
rect 45928 9036 45980 9042
rect 45928 8978 45980 8984
rect 46020 9036 46072 9042
rect 46020 8978 46072 8984
rect 46112 8968 46164 8974
rect 46018 8936 46074 8945
rect 46112 8910 46164 8916
rect 46018 8871 46074 8880
rect 46032 8498 46060 8871
rect 46124 8634 46152 8910
rect 46216 8906 46244 9454
rect 46294 9415 46350 9424
rect 46400 9178 46428 12135
rect 46492 10538 46520 16526
rect 46584 12345 46612 17190
rect 46848 16584 46900 16590
rect 46848 16526 46900 16532
rect 46756 16516 46808 16522
rect 46756 16458 46808 16464
rect 46664 16040 46716 16046
rect 46664 15982 46716 15988
rect 46676 15570 46704 15982
rect 46768 15978 46796 16458
rect 46860 16114 46888 16526
rect 46848 16108 46900 16114
rect 46848 16050 46900 16056
rect 46756 15972 46808 15978
rect 46756 15914 46808 15920
rect 46846 15600 46902 15609
rect 46664 15564 46716 15570
rect 46846 15535 46902 15544
rect 46664 15506 46716 15512
rect 46676 15348 46704 15506
rect 46860 15502 46888 15535
rect 46848 15496 46900 15502
rect 46848 15438 46900 15444
rect 46756 15360 46808 15366
rect 46676 15320 46756 15348
rect 46756 15302 46808 15308
rect 46664 14952 46716 14958
rect 46662 14920 46664 14929
rect 46716 14920 46718 14929
rect 46662 14855 46718 14864
rect 46664 14476 46716 14482
rect 46664 14418 46716 14424
rect 46676 14385 46704 14418
rect 46662 14376 46718 14385
rect 46662 14311 46718 14320
rect 46664 13932 46716 13938
rect 46664 13874 46716 13880
rect 46676 13841 46704 13874
rect 46768 13870 46796 15302
rect 46846 15192 46902 15201
rect 46846 15127 46902 15136
rect 46860 14074 46888 15127
rect 46952 14618 46980 18702
rect 47216 18624 47268 18630
rect 47216 18566 47268 18572
rect 47124 17332 47176 17338
rect 47124 17274 47176 17280
rect 47032 16040 47084 16046
rect 47032 15982 47084 15988
rect 47044 15502 47072 15982
rect 47032 15496 47084 15502
rect 47032 15438 47084 15444
rect 47032 14816 47084 14822
rect 47032 14758 47084 14764
rect 46940 14612 46992 14618
rect 46940 14554 46992 14560
rect 47044 14414 47072 14758
rect 47136 14414 47164 17274
rect 47228 17134 47256 18566
rect 47320 17762 47348 22646
rect 47596 22094 47624 26318
rect 48056 26314 48176 26330
rect 48780 26376 48832 26382
rect 48780 26318 48832 26324
rect 49148 26376 49200 26382
rect 49148 26318 49200 26324
rect 49240 26376 49292 26382
rect 49240 26318 49292 26324
rect 49516 26376 49568 26382
rect 49516 26318 49568 26324
rect 50620 26376 50672 26382
rect 50620 26318 50672 26324
rect 50712 26376 50764 26382
rect 50712 26318 50764 26324
rect 48044 26308 48176 26314
rect 48096 26302 48176 26308
rect 48044 26250 48096 26256
rect 48056 26042 48084 26250
rect 48792 26058 48820 26318
rect 48044 26036 48096 26042
rect 48792 26030 48912 26058
rect 48044 25978 48096 25984
rect 48780 25968 48832 25974
rect 48780 25910 48832 25916
rect 47676 25696 47728 25702
rect 47676 25638 47728 25644
rect 47688 22438 47716 25638
rect 48792 25498 48820 25910
rect 48884 25906 48912 26030
rect 48872 25900 48924 25906
rect 48872 25842 48924 25848
rect 49160 25702 49188 26318
rect 49252 25838 49280 26318
rect 49424 25900 49476 25906
rect 49424 25842 49476 25848
rect 49240 25832 49292 25838
rect 49240 25774 49292 25780
rect 49148 25696 49200 25702
rect 49148 25638 49200 25644
rect 48780 25492 48832 25498
rect 48780 25434 48832 25440
rect 48504 25288 48556 25294
rect 48504 25230 48556 25236
rect 48516 24954 48544 25230
rect 48964 25220 49016 25226
rect 48964 25162 49016 25168
rect 48504 24948 48556 24954
rect 48504 24890 48556 24896
rect 48516 24857 48544 24890
rect 48502 24848 48558 24857
rect 48502 24783 48558 24792
rect 48976 24614 49004 25162
rect 48964 24608 49016 24614
rect 48964 24550 49016 24556
rect 48596 23792 48648 23798
rect 48596 23734 48648 23740
rect 48964 23792 49016 23798
rect 48964 23734 49016 23740
rect 48608 23662 48636 23734
rect 48596 23656 48648 23662
rect 48596 23598 48648 23604
rect 48044 23180 48096 23186
rect 48044 23122 48096 23128
rect 48056 22778 48084 23122
rect 48608 22982 48636 23598
rect 48688 23520 48740 23526
rect 48688 23462 48740 23468
rect 48700 23118 48728 23462
rect 48976 23118 49004 23734
rect 49160 23322 49188 25638
rect 49252 23526 49280 25774
rect 49436 24954 49464 25842
rect 49528 25770 49556 26318
rect 50816 26314 50844 26982
rect 51000 26586 51028 27798
rect 51184 27130 51212 27968
rect 51368 27674 51396 28018
rect 51356 27668 51408 27674
rect 51356 27610 51408 27616
rect 52932 27538 52960 28036
rect 53012 28076 53064 28082
rect 53012 28018 53064 28024
rect 53748 28076 53800 28082
rect 53748 28018 53800 28024
rect 52276 27532 52328 27538
rect 52276 27474 52328 27480
rect 52920 27532 52972 27538
rect 52920 27474 52972 27480
rect 51172 27124 51224 27130
rect 51172 27066 51224 27072
rect 52288 26994 52316 27474
rect 52368 27464 52420 27470
rect 52368 27406 52420 27412
rect 52380 26994 52408 27406
rect 53024 27062 53052 28018
rect 53196 27872 53248 27878
rect 53196 27814 53248 27820
rect 53012 27056 53064 27062
rect 53012 26998 53064 27004
rect 52276 26988 52328 26994
rect 52276 26930 52328 26936
rect 52368 26988 52420 26994
rect 52368 26930 52420 26936
rect 50988 26580 51040 26586
rect 50988 26522 51040 26528
rect 49608 26308 49660 26314
rect 49608 26250 49660 26256
rect 50804 26308 50856 26314
rect 50804 26250 50856 26256
rect 49620 25974 49648 26250
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 49608 25968 49660 25974
rect 49608 25910 49660 25916
rect 49884 25900 49936 25906
rect 49884 25842 49936 25848
rect 50712 25900 50764 25906
rect 50712 25842 50764 25848
rect 49516 25764 49568 25770
rect 49516 25706 49568 25712
rect 49516 25288 49568 25294
rect 49516 25230 49568 25236
rect 49424 24948 49476 24954
rect 49424 24890 49476 24896
rect 49528 24818 49556 25230
rect 49792 25152 49844 25158
rect 49792 25094 49844 25100
rect 49804 24886 49832 25094
rect 49792 24880 49844 24886
rect 49792 24822 49844 24828
rect 49516 24812 49568 24818
rect 49516 24754 49568 24760
rect 49804 23746 49832 24822
rect 49896 24818 49924 25842
rect 50724 25362 50752 25842
rect 50816 25498 50844 26250
rect 52288 26234 52316 26930
rect 52196 26206 52316 26234
rect 50988 25900 51040 25906
rect 50988 25842 51040 25848
rect 50804 25492 50856 25498
rect 50804 25434 50856 25440
rect 50712 25356 50764 25362
rect 50712 25298 50764 25304
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 49884 24812 49936 24818
rect 49884 24754 49936 24760
rect 49896 23866 49924 24754
rect 49976 24744 50028 24750
rect 49976 24686 50028 24692
rect 49884 23860 49936 23866
rect 49884 23802 49936 23808
rect 49700 23724 49752 23730
rect 49804 23718 49924 23746
rect 49988 23730 50016 24686
rect 50068 24676 50120 24682
rect 50068 24618 50120 24624
rect 50080 23798 50108 24618
rect 50160 24608 50212 24614
rect 50160 24550 50212 24556
rect 50068 23792 50120 23798
rect 50068 23734 50120 23740
rect 49700 23666 49752 23672
rect 49424 23656 49476 23662
rect 49424 23598 49476 23604
rect 49240 23520 49292 23526
rect 49240 23462 49292 23468
rect 49148 23316 49200 23322
rect 49148 23258 49200 23264
rect 48688 23112 48740 23118
rect 48688 23054 48740 23060
rect 48964 23112 49016 23118
rect 48964 23054 49016 23060
rect 48596 22976 48648 22982
rect 48596 22918 48648 22924
rect 48044 22772 48096 22778
rect 48044 22714 48096 22720
rect 47676 22432 47728 22438
rect 47676 22374 47728 22380
rect 47504 22066 47624 22094
rect 47504 21078 47532 22066
rect 47492 21072 47544 21078
rect 47492 21014 47544 21020
rect 47400 20868 47452 20874
rect 47400 20810 47452 20816
rect 47412 20058 47440 20810
rect 47400 20052 47452 20058
rect 47400 19994 47452 20000
rect 47492 19780 47544 19786
rect 47492 19722 47544 19728
rect 47504 18970 47532 19722
rect 47492 18964 47544 18970
rect 47492 18906 47544 18912
rect 47584 18760 47636 18766
rect 47584 18702 47636 18708
rect 47596 18154 47624 18702
rect 47584 18148 47636 18154
rect 47584 18090 47636 18096
rect 47492 17876 47544 17882
rect 47492 17818 47544 17824
rect 47320 17734 47440 17762
rect 47308 17672 47360 17678
rect 47308 17614 47360 17620
rect 47216 17128 47268 17134
rect 47216 17070 47268 17076
rect 47228 16289 47256 17070
rect 47214 16280 47270 16289
rect 47214 16215 47216 16224
rect 47268 16215 47270 16224
rect 47216 16186 47268 16192
rect 47228 16155 47256 16186
rect 47320 16153 47348 17614
rect 47412 17610 47440 17734
rect 47400 17604 47452 17610
rect 47400 17546 47452 17552
rect 47398 16688 47454 16697
rect 47398 16623 47454 16632
rect 47412 16590 47440 16623
rect 47400 16584 47452 16590
rect 47400 16526 47452 16532
rect 47306 16144 47362 16153
rect 47306 16079 47362 16088
rect 47400 16108 47452 16114
rect 47400 16050 47452 16056
rect 47412 15706 47440 16050
rect 47400 15700 47452 15706
rect 47400 15642 47452 15648
rect 47412 15570 47440 15642
rect 47504 15570 47532 17818
rect 47582 17640 47638 17649
rect 47582 17575 47638 17584
rect 47596 17542 47624 17575
rect 47584 17536 47636 17542
rect 47584 17478 47636 17484
rect 47400 15564 47452 15570
rect 47320 15524 47400 15552
rect 47216 14816 47268 14822
rect 47216 14758 47268 14764
rect 47032 14408 47084 14414
rect 47032 14350 47084 14356
rect 47124 14408 47176 14414
rect 47124 14350 47176 14356
rect 46940 14340 46992 14346
rect 46940 14282 46992 14288
rect 46848 14068 46900 14074
rect 46848 14010 46900 14016
rect 46860 13938 46888 14010
rect 46848 13932 46900 13938
rect 46848 13874 46900 13880
rect 46756 13864 46808 13870
rect 46662 13832 46718 13841
rect 46756 13806 46808 13812
rect 46662 13767 46718 13776
rect 46676 12782 46704 13767
rect 46768 13394 46796 13806
rect 46756 13388 46808 13394
rect 46756 13330 46808 13336
rect 46754 13152 46810 13161
rect 46754 13087 46810 13096
rect 46768 12782 46796 13087
rect 46664 12776 46716 12782
rect 46664 12718 46716 12724
rect 46756 12776 46808 12782
rect 46756 12718 46808 12724
rect 46664 12640 46716 12646
rect 46664 12582 46716 12588
rect 46570 12336 46626 12345
rect 46570 12271 46626 12280
rect 46676 12170 46704 12582
rect 46664 12164 46716 12170
rect 46664 12106 46716 12112
rect 46768 11676 46796 12718
rect 46848 12164 46900 12170
rect 46848 12106 46900 12112
rect 46860 11898 46888 12106
rect 46848 11892 46900 11898
rect 46848 11834 46900 11840
rect 46676 11648 46796 11676
rect 46676 10674 46704 11648
rect 46756 11552 46808 11558
rect 46756 11494 46808 11500
rect 46664 10668 46716 10674
rect 46664 10610 46716 10616
rect 46572 10600 46624 10606
rect 46572 10542 46624 10548
rect 46480 10532 46532 10538
rect 46480 10474 46532 10480
rect 46480 9716 46532 9722
rect 46480 9658 46532 9664
rect 46492 9450 46520 9658
rect 46480 9444 46532 9450
rect 46480 9386 46532 9392
rect 46388 9172 46440 9178
rect 46388 9114 46440 9120
rect 46294 9072 46350 9081
rect 46294 9007 46350 9016
rect 46308 8974 46336 9007
rect 46296 8968 46348 8974
rect 46296 8910 46348 8916
rect 46204 8900 46256 8906
rect 46204 8842 46256 8848
rect 46112 8628 46164 8634
rect 46112 8570 46164 8576
rect 46216 8566 46244 8842
rect 46204 8560 46256 8566
rect 46204 8502 46256 8508
rect 46020 8492 46072 8498
rect 46020 8434 46072 8440
rect 46492 8090 46520 9386
rect 46584 8838 46612 10542
rect 46664 10532 46716 10538
rect 46664 10474 46716 10480
rect 46572 8832 46624 8838
rect 46572 8774 46624 8780
rect 46572 8560 46624 8566
rect 46572 8502 46624 8508
rect 46584 8362 46612 8502
rect 46676 8498 46704 10474
rect 46768 10130 46796 11494
rect 46952 11354 46980 14282
rect 47032 14068 47084 14074
rect 47032 14010 47084 14016
rect 47044 13258 47072 14010
rect 47136 13530 47164 14350
rect 47124 13524 47176 13530
rect 47124 13466 47176 13472
rect 47228 13462 47256 14758
rect 47216 13456 47268 13462
rect 47216 13398 47268 13404
rect 47032 13252 47084 13258
rect 47032 13194 47084 13200
rect 47044 13161 47072 13194
rect 47030 13152 47086 13161
rect 47030 13087 47086 13096
rect 47320 12986 47348 15524
rect 47400 15506 47452 15512
rect 47492 15564 47544 15570
rect 47492 15506 47544 15512
rect 47400 15428 47452 15434
rect 47400 15370 47452 15376
rect 47412 15094 47440 15370
rect 47400 15088 47452 15094
rect 47400 15030 47452 15036
rect 47400 14408 47452 14414
rect 47400 14350 47452 14356
rect 47412 14074 47440 14350
rect 47400 14068 47452 14074
rect 47400 14010 47452 14016
rect 47400 13932 47452 13938
rect 47400 13874 47452 13880
rect 47412 13705 47440 13874
rect 47398 13696 47454 13705
rect 47398 13631 47454 13640
rect 47308 12980 47360 12986
rect 47308 12922 47360 12928
rect 47216 12844 47268 12850
rect 47216 12786 47268 12792
rect 47032 12232 47084 12238
rect 47032 12174 47084 12180
rect 46940 11348 46992 11354
rect 46940 11290 46992 11296
rect 46848 10804 46900 10810
rect 46952 10792 46980 11290
rect 46900 10764 46980 10792
rect 46848 10746 46900 10752
rect 47044 10538 47072 12174
rect 47124 12164 47176 12170
rect 47124 12106 47176 12112
rect 47032 10532 47084 10538
rect 47032 10474 47084 10480
rect 46940 10464 46992 10470
rect 46940 10406 46992 10412
rect 46846 10160 46902 10169
rect 46756 10124 46808 10130
rect 46846 10095 46902 10104
rect 46756 10066 46808 10072
rect 46860 10062 46888 10095
rect 46848 10056 46900 10062
rect 46848 9998 46900 10004
rect 46756 9988 46808 9994
rect 46756 9930 46808 9936
rect 46664 8492 46716 8498
rect 46664 8434 46716 8440
rect 46572 8356 46624 8362
rect 46572 8298 46624 8304
rect 46480 8084 46532 8090
rect 46480 8026 46532 8032
rect 46572 8084 46624 8090
rect 46572 8026 46624 8032
rect 46388 8016 46440 8022
rect 46388 7958 46440 7964
rect 45836 7744 45888 7750
rect 45836 7686 45888 7692
rect 46296 7744 46348 7750
rect 46296 7686 46348 7692
rect 45744 7540 45796 7546
rect 45744 7482 45796 7488
rect 45744 6996 45796 7002
rect 45744 6938 45796 6944
rect 45756 6730 45784 6938
rect 45744 6724 45796 6730
rect 45744 6666 45796 6672
rect 45652 5636 45704 5642
rect 45652 5578 45704 5584
rect 45560 5296 45612 5302
rect 45560 5238 45612 5244
rect 45480 5086 45600 5114
rect 45572 4010 45600 5086
rect 45664 4486 45692 5578
rect 45756 5574 45784 6666
rect 45744 5568 45796 5574
rect 45744 5510 45796 5516
rect 45848 5166 45876 7686
rect 46308 7478 46336 7686
rect 46400 7478 46428 7958
rect 46584 7886 46612 8026
rect 46572 7880 46624 7886
rect 46572 7822 46624 7828
rect 46480 7744 46532 7750
rect 46480 7686 46532 7692
rect 46296 7472 46348 7478
rect 46296 7414 46348 7420
rect 46388 7472 46440 7478
rect 46388 7414 46440 7420
rect 46204 7404 46256 7410
rect 46204 7346 46256 7352
rect 45928 6656 45980 6662
rect 45928 6598 45980 6604
rect 45940 6118 45968 6598
rect 45928 6112 45980 6118
rect 45928 6054 45980 6060
rect 46216 5914 46244 7346
rect 46388 7336 46440 7342
rect 46492 7324 46520 7686
rect 46440 7296 46520 7324
rect 46388 7278 46440 7284
rect 46296 6656 46348 6662
rect 46296 6598 46348 6604
rect 46308 6322 46336 6598
rect 46296 6316 46348 6322
rect 46296 6258 46348 6264
rect 46388 6316 46440 6322
rect 46388 6258 46440 6264
rect 46204 5908 46256 5914
rect 46204 5850 46256 5856
rect 46400 5778 46428 6258
rect 46388 5772 46440 5778
rect 46388 5714 46440 5720
rect 46018 5672 46074 5681
rect 46018 5607 46074 5616
rect 46032 5574 46060 5607
rect 46020 5568 46072 5574
rect 46020 5510 46072 5516
rect 45836 5160 45888 5166
rect 45836 5102 45888 5108
rect 45848 4826 45876 5102
rect 45744 4820 45796 4826
rect 45744 4762 45796 4768
rect 45836 4820 45888 4826
rect 45836 4762 45888 4768
rect 45756 4690 45784 4762
rect 45744 4684 45796 4690
rect 45744 4626 45796 4632
rect 45652 4480 45704 4486
rect 45652 4422 45704 4428
rect 45756 4146 45784 4626
rect 45744 4140 45796 4146
rect 45744 4082 45796 4088
rect 45560 4004 45612 4010
rect 45560 3946 45612 3952
rect 45652 3936 45704 3942
rect 45652 3878 45704 3884
rect 45284 3120 45336 3126
rect 45284 3062 45336 3068
rect 45376 3120 45428 3126
rect 45376 3062 45428 3068
rect 45192 2644 45244 2650
rect 45192 2586 45244 2592
rect 45664 2582 45692 3878
rect 45848 3754 45876 4762
rect 46032 4554 46060 5510
rect 46386 5128 46442 5137
rect 46386 5063 46442 5072
rect 46204 5024 46256 5030
rect 46204 4966 46256 4972
rect 46020 4548 46072 4554
rect 46020 4490 46072 4496
rect 45928 4480 45980 4486
rect 45928 4422 45980 4428
rect 45756 3726 45876 3754
rect 45756 3670 45784 3726
rect 45744 3664 45796 3670
rect 45744 3606 45796 3612
rect 45940 3398 45968 4422
rect 46216 4282 46244 4966
rect 46400 4486 46428 5063
rect 46492 5030 46520 7296
rect 46676 6934 46704 8434
rect 46768 7954 46796 9930
rect 46848 9580 46900 9586
rect 46848 9522 46900 9528
rect 46860 8498 46888 9522
rect 46952 9382 46980 10406
rect 47136 9654 47164 12106
rect 47228 11937 47256 12786
rect 47214 11928 47270 11937
rect 47214 11863 47270 11872
rect 47216 11824 47268 11830
rect 47216 11766 47268 11772
rect 47228 11286 47256 11766
rect 47216 11280 47268 11286
rect 47216 11222 47268 11228
rect 47320 11150 47348 12922
rect 47412 11898 47440 13631
rect 47400 11892 47452 11898
rect 47400 11834 47452 11840
rect 47504 11218 47532 15506
rect 47596 15502 47624 17478
rect 47584 15496 47636 15502
rect 47584 15438 47636 15444
rect 47492 11212 47544 11218
rect 47492 11154 47544 11160
rect 47308 11144 47360 11150
rect 47308 11086 47360 11092
rect 47400 11076 47452 11082
rect 47400 11018 47452 11024
rect 47124 9648 47176 9654
rect 47124 9590 47176 9596
rect 46940 9376 46992 9382
rect 46940 9318 46992 9324
rect 46848 8492 46900 8498
rect 46848 8434 46900 8440
rect 46952 8294 46980 9318
rect 47032 9104 47084 9110
rect 47030 9072 47032 9081
rect 47084 9072 47086 9081
rect 47030 9007 47086 9016
rect 47136 8362 47164 9590
rect 47412 9353 47440 11018
rect 47398 9344 47454 9353
rect 47398 9279 47454 9288
rect 47216 8968 47268 8974
rect 47216 8910 47268 8916
rect 47306 8936 47362 8945
rect 47124 8356 47176 8362
rect 47124 8298 47176 8304
rect 46940 8288 46992 8294
rect 47228 8242 47256 8910
rect 47306 8871 47362 8880
rect 46940 8230 46992 8236
rect 47136 8214 47256 8242
rect 46756 7948 46808 7954
rect 46756 7890 46808 7896
rect 46768 7313 46796 7890
rect 46940 7472 46992 7478
rect 46940 7414 46992 7420
rect 46754 7304 46810 7313
rect 46754 7239 46810 7248
rect 46952 7002 46980 7414
rect 47032 7200 47084 7206
rect 47032 7142 47084 7148
rect 46940 6996 46992 7002
rect 46940 6938 46992 6944
rect 46572 6928 46624 6934
rect 46572 6870 46624 6876
rect 46664 6928 46716 6934
rect 46664 6870 46716 6876
rect 46584 5273 46612 6870
rect 46756 6860 46808 6866
rect 46756 6802 46808 6808
rect 46768 6322 46796 6802
rect 46848 6384 46900 6390
rect 46848 6326 46900 6332
rect 46756 6316 46808 6322
rect 46756 6258 46808 6264
rect 46860 5370 46888 6326
rect 47044 6322 47072 7142
rect 47032 6316 47084 6322
rect 47032 6258 47084 6264
rect 46940 5568 46992 5574
rect 47136 5556 47164 8214
rect 47216 7404 47268 7410
rect 47216 7346 47268 7352
rect 47228 7002 47256 7346
rect 47216 6996 47268 7002
rect 47216 6938 47268 6944
rect 47320 6798 47348 8871
rect 47400 6860 47452 6866
rect 47400 6802 47452 6808
rect 47308 6792 47360 6798
rect 47308 6734 47360 6740
rect 47320 6186 47348 6734
rect 47412 6662 47440 6802
rect 47400 6656 47452 6662
rect 47400 6598 47452 6604
rect 47308 6180 47360 6186
rect 47308 6122 47360 6128
rect 47216 5704 47268 5710
rect 47320 5692 47348 6122
rect 47268 5664 47348 5692
rect 47216 5646 47268 5652
rect 47504 5642 47532 11154
rect 47596 11150 47624 15438
rect 47584 11144 47636 11150
rect 47584 11086 47636 11092
rect 47596 8945 47624 11086
rect 47688 10266 47716 22374
rect 48976 22234 49004 23054
rect 49436 23050 49464 23598
rect 49712 23254 49740 23666
rect 49792 23520 49844 23526
rect 49792 23462 49844 23468
rect 49700 23248 49752 23254
rect 49700 23190 49752 23196
rect 49804 23118 49832 23462
rect 49792 23112 49844 23118
rect 49792 23054 49844 23060
rect 49424 23044 49476 23050
rect 49424 22986 49476 22992
rect 49240 22636 49292 22642
rect 49240 22578 49292 22584
rect 48964 22228 49016 22234
rect 48964 22170 49016 22176
rect 49252 22098 49280 22578
rect 49436 22438 49464 22986
rect 49700 22568 49752 22574
rect 49700 22510 49752 22516
rect 49424 22432 49476 22438
rect 49424 22374 49476 22380
rect 49436 22098 49464 22374
rect 47768 22092 47820 22098
rect 47768 22034 47820 22040
rect 47860 22092 47912 22098
rect 47860 22034 47912 22040
rect 49240 22092 49292 22098
rect 49240 22034 49292 22040
rect 49424 22092 49476 22098
rect 49424 22034 49476 22040
rect 47780 21690 47808 22034
rect 47768 21684 47820 21690
rect 47768 21626 47820 21632
rect 47872 21554 47900 22034
rect 48780 22024 48832 22030
rect 48780 21966 48832 21972
rect 49148 22024 49200 22030
rect 49148 21966 49200 21972
rect 48792 21690 48820 21966
rect 48780 21684 48832 21690
rect 48780 21626 48832 21632
rect 47768 21548 47820 21554
rect 47768 21490 47820 21496
rect 47860 21548 47912 21554
rect 47860 21490 47912 21496
rect 48228 21548 48280 21554
rect 48228 21490 48280 21496
rect 47780 19990 47808 21490
rect 47768 19984 47820 19990
rect 47768 19926 47820 19932
rect 47872 19718 47900 21490
rect 48240 20942 48268 21490
rect 48964 21344 49016 21350
rect 48964 21286 49016 21292
rect 48976 20942 49004 21286
rect 49160 21146 49188 21966
rect 49252 21690 49280 22034
rect 49240 21684 49292 21690
rect 49240 21626 49292 21632
rect 49240 21548 49292 21554
rect 49240 21490 49292 21496
rect 49148 21140 49200 21146
rect 49148 21082 49200 21088
rect 47952 20936 48004 20942
rect 47952 20878 48004 20884
rect 48136 20936 48188 20942
rect 48136 20878 48188 20884
rect 48228 20936 48280 20942
rect 48228 20878 48280 20884
rect 48964 20936 49016 20942
rect 49148 20936 49200 20942
rect 48964 20878 49016 20884
rect 49146 20904 49148 20913
rect 49252 20924 49280 21490
rect 49200 20904 49280 20924
rect 49202 20896 49280 20904
rect 47964 20534 47992 20878
rect 47952 20528 48004 20534
rect 47952 20470 48004 20476
rect 48148 20466 48176 20878
rect 48976 20602 49004 20878
rect 49146 20839 49202 20848
rect 48964 20596 49016 20602
rect 48964 20538 49016 20544
rect 48136 20460 48188 20466
rect 48136 20402 48188 20408
rect 48780 20460 48832 20466
rect 48780 20402 48832 20408
rect 47860 19712 47912 19718
rect 47860 19654 47912 19660
rect 48148 19310 48176 20402
rect 48596 19984 48648 19990
rect 48596 19926 48648 19932
rect 48228 19848 48280 19854
rect 48228 19790 48280 19796
rect 48240 19514 48268 19790
rect 48608 19786 48636 19926
rect 48596 19780 48648 19786
rect 48596 19722 48648 19728
rect 48608 19514 48636 19722
rect 48228 19508 48280 19514
rect 48228 19450 48280 19456
rect 48596 19508 48648 19514
rect 48596 19450 48648 19456
rect 48136 19304 48188 19310
rect 47964 19264 48136 19292
rect 47964 17954 47992 19264
rect 48136 19246 48188 19252
rect 48504 18284 48556 18290
rect 48504 18226 48556 18232
rect 48412 18080 48464 18086
rect 48412 18022 48464 18028
rect 47964 17926 48084 17954
rect 47768 17808 47820 17814
rect 47768 17750 47820 17756
rect 47780 17678 47808 17750
rect 47768 17672 47820 17678
rect 47768 17614 47820 17620
rect 47860 16788 47912 16794
rect 47860 16730 47912 16736
rect 47872 16590 47900 16730
rect 48056 16726 48084 17926
rect 48320 17604 48372 17610
rect 48320 17546 48372 17552
rect 48332 17270 48360 17546
rect 48320 17264 48372 17270
rect 48320 17206 48372 17212
rect 48318 17096 48374 17105
rect 48318 17031 48320 17040
rect 48372 17031 48374 17040
rect 48320 17002 48372 17008
rect 48424 16726 48452 18022
rect 48516 17882 48544 18226
rect 48504 17876 48556 17882
rect 48504 17818 48556 17824
rect 48504 17128 48556 17134
rect 48502 17096 48504 17105
rect 48556 17096 48558 17105
rect 48502 17031 48558 17040
rect 48044 16720 48096 16726
rect 48044 16662 48096 16668
rect 48412 16720 48464 16726
rect 48412 16662 48464 16668
rect 47860 16584 47912 16590
rect 47860 16526 47912 16532
rect 48274 16448 48326 16454
rect 48504 16448 48556 16454
rect 48326 16396 48452 16402
rect 48274 16390 48452 16396
rect 48504 16390 48556 16396
rect 48286 16374 48452 16390
rect 48318 16280 48374 16289
rect 48318 16215 48374 16224
rect 47860 16176 47912 16182
rect 47860 16118 47912 16124
rect 47872 15609 47900 16118
rect 48136 16108 48188 16114
rect 48136 16050 48188 16056
rect 47952 15972 48004 15978
rect 47952 15914 48004 15920
rect 47964 15881 47992 15914
rect 47950 15872 48006 15881
rect 47950 15807 48006 15816
rect 47952 15632 48004 15638
rect 47858 15600 47914 15609
rect 47768 15564 47820 15570
rect 47952 15574 48004 15580
rect 47858 15535 47914 15544
rect 47768 15506 47820 15512
rect 47780 15201 47808 15506
rect 47860 15360 47912 15366
rect 47860 15302 47912 15308
rect 47766 15192 47822 15201
rect 47872 15162 47900 15302
rect 47766 15127 47822 15136
rect 47860 15156 47912 15162
rect 47860 15098 47912 15104
rect 47768 15088 47820 15094
rect 47768 15030 47820 15036
rect 47780 14346 47808 15030
rect 47768 14340 47820 14346
rect 47768 14282 47820 14288
rect 47860 14068 47912 14074
rect 47860 14010 47912 14016
rect 47768 13864 47820 13870
rect 47768 13806 47820 13812
rect 47780 11830 47808 13806
rect 47872 13161 47900 14010
rect 47964 13394 47992 15574
rect 48044 15020 48096 15026
rect 48044 14962 48096 14968
rect 48056 14618 48084 14962
rect 48044 14612 48096 14618
rect 48044 14554 48096 14560
rect 48042 13560 48098 13569
rect 48042 13495 48044 13504
rect 48096 13495 48098 13504
rect 48044 13466 48096 13472
rect 47952 13388 48004 13394
rect 47952 13330 48004 13336
rect 48148 13326 48176 16050
rect 48228 15496 48280 15502
rect 48228 15438 48280 15444
rect 48240 14822 48268 15438
rect 48228 14816 48280 14822
rect 48228 14758 48280 14764
rect 48332 14346 48360 16215
rect 48424 15745 48452 16374
rect 48516 16250 48544 16390
rect 48504 16244 48556 16250
rect 48504 16186 48556 16192
rect 48502 15872 48558 15881
rect 48502 15807 48558 15816
rect 48410 15736 48466 15745
rect 48410 15671 48466 15680
rect 48516 15162 48544 15807
rect 48504 15156 48556 15162
rect 48504 15098 48556 15104
rect 48412 14884 48464 14890
rect 48412 14826 48464 14832
rect 48504 14884 48556 14890
rect 48504 14826 48556 14832
rect 48424 14414 48452 14826
rect 48516 14793 48544 14826
rect 48502 14784 48558 14793
rect 48502 14719 48558 14728
rect 48412 14408 48464 14414
rect 48412 14350 48464 14356
rect 48502 14376 48558 14385
rect 48320 14340 48372 14346
rect 48502 14311 48558 14320
rect 48320 14282 48372 14288
rect 48226 13696 48282 13705
rect 48226 13631 48282 13640
rect 48240 13326 48268 13631
rect 48136 13320 48188 13326
rect 48136 13262 48188 13268
rect 48228 13320 48280 13326
rect 48228 13262 48280 13268
rect 48044 13252 48096 13258
rect 48044 13194 48096 13200
rect 47858 13152 47914 13161
rect 47858 13087 47914 13096
rect 48056 12850 48084 13194
rect 48044 12844 48096 12850
rect 48044 12786 48096 12792
rect 48056 12434 48084 12786
rect 48148 12646 48176 13262
rect 48228 12912 48280 12918
rect 48228 12854 48280 12860
rect 48136 12640 48188 12646
rect 48136 12582 48188 12588
rect 47872 12406 48084 12434
rect 48136 12436 48188 12442
rect 47768 11824 47820 11830
rect 47768 11766 47820 11772
rect 47768 11348 47820 11354
rect 47768 11290 47820 11296
rect 47780 11150 47808 11290
rect 47768 11144 47820 11150
rect 47768 11086 47820 11092
rect 47780 10674 47808 11086
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 47872 10554 47900 12406
rect 48136 12378 48188 12384
rect 48148 12306 48176 12378
rect 48136 12300 48188 12306
rect 48136 12242 48188 12248
rect 48044 11008 48096 11014
rect 48044 10950 48096 10956
rect 48056 10742 48084 10950
rect 48044 10736 48096 10742
rect 48044 10678 48096 10684
rect 47780 10526 47900 10554
rect 47676 10260 47728 10266
rect 47676 10202 47728 10208
rect 47582 8936 47638 8945
rect 47582 8871 47638 8880
rect 47780 8838 47808 10526
rect 48148 10062 48176 12242
rect 48240 12102 48268 12854
rect 48332 12850 48360 14282
rect 48516 14260 48544 14311
rect 48424 14232 48544 14260
rect 48424 13734 48452 14232
rect 48504 13932 48556 13938
rect 48504 13874 48556 13880
rect 48412 13728 48464 13734
rect 48412 13670 48464 13676
rect 48424 12918 48452 13670
rect 48516 13569 48544 13874
rect 48502 13560 48558 13569
rect 48502 13495 48504 13504
rect 48556 13495 48558 13504
rect 48504 13466 48556 13472
rect 48608 13410 48636 19450
rect 48792 19242 48820 20402
rect 48872 20324 48924 20330
rect 48872 20266 48924 20272
rect 48884 19854 48912 20266
rect 48976 19922 49004 20538
rect 49148 20256 49200 20262
rect 49148 20198 49200 20204
rect 49160 20058 49188 20198
rect 49148 20052 49200 20058
rect 49148 19994 49200 20000
rect 48964 19916 49016 19922
rect 48964 19858 49016 19864
rect 48872 19848 48924 19854
rect 48872 19790 48924 19796
rect 49148 19780 49200 19786
rect 49148 19722 49200 19728
rect 49160 19242 49188 19722
rect 48780 19236 48832 19242
rect 48780 19178 48832 19184
rect 49148 19236 49200 19242
rect 49148 19178 49200 19184
rect 48964 18284 49016 18290
rect 48964 18226 49016 18232
rect 48976 17814 49004 18226
rect 48964 17808 49016 17814
rect 48964 17750 49016 17756
rect 48872 17536 48924 17542
rect 48872 17478 48924 17484
rect 48884 17202 48912 17478
rect 48872 17196 48924 17202
rect 48872 17138 48924 17144
rect 48964 17196 49016 17202
rect 48964 17138 49016 17144
rect 48778 16688 48834 16697
rect 48976 16640 49004 17138
rect 49056 17128 49108 17134
rect 49056 17070 49108 17076
rect 48778 16623 48780 16632
rect 48832 16623 48834 16632
rect 48780 16594 48832 16600
rect 48884 16612 49004 16640
rect 48780 16516 48832 16522
rect 48780 16458 48832 16464
rect 48688 16108 48740 16114
rect 48688 16050 48740 16056
rect 48700 15706 48728 16050
rect 48792 15881 48820 16458
rect 48778 15872 48834 15881
rect 48778 15807 48834 15816
rect 48688 15700 48740 15706
rect 48688 15642 48740 15648
rect 48884 15484 48912 16612
rect 48962 16280 49018 16289
rect 48962 16215 49018 16224
rect 48976 16046 49004 16215
rect 48964 16040 49016 16046
rect 48964 15982 49016 15988
rect 48964 15904 49016 15910
rect 48964 15846 49016 15852
rect 48700 15456 48912 15484
rect 48700 14958 48728 15456
rect 48780 15020 48832 15026
rect 48780 14962 48832 14968
rect 48688 14952 48740 14958
rect 48688 14894 48740 14900
rect 48700 14550 48728 14894
rect 48792 14793 48820 14962
rect 48872 14952 48924 14958
rect 48872 14894 48924 14900
rect 48778 14784 48834 14793
rect 48778 14719 48834 14728
rect 48688 14544 48740 14550
rect 48688 14486 48740 14492
rect 48688 14408 48740 14414
rect 48688 14350 48740 14356
rect 48700 13530 48728 14350
rect 48792 13852 48820 14719
rect 48884 14618 48912 14894
rect 48872 14612 48924 14618
rect 48872 14554 48924 14560
rect 48976 14385 49004 15846
rect 49068 14414 49096 17070
rect 49056 14408 49108 14414
rect 48962 14376 49018 14385
rect 49056 14350 49108 14356
rect 48962 14311 49018 14320
rect 49056 14272 49108 14278
rect 49056 14214 49108 14220
rect 48792 13824 48912 13852
rect 48688 13524 48740 13530
rect 48688 13466 48740 13472
rect 48504 13388 48556 13394
rect 48608 13382 48820 13410
rect 48504 13330 48556 13336
rect 48516 13258 48544 13330
rect 48594 13288 48650 13297
rect 48504 13252 48556 13258
rect 48594 13223 48650 13232
rect 48688 13252 48740 13258
rect 48504 13194 48556 13200
rect 48412 12912 48464 12918
rect 48412 12854 48464 12860
rect 48320 12844 48372 12850
rect 48320 12786 48372 12792
rect 48318 12472 48374 12481
rect 48608 12442 48636 13223
rect 48688 13194 48740 13200
rect 48318 12407 48374 12416
rect 48596 12436 48648 12442
rect 48332 12374 48360 12407
rect 48596 12378 48648 12384
rect 48320 12368 48372 12374
rect 48504 12368 48556 12374
rect 48320 12310 48372 12316
rect 48410 12336 48466 12345
rect 48504 12310 48556 12316
rect 48700 12322 48728 13194
rect 48792 12442 48820 13382
rect 48780 12436 48832 12442
rect 48780 12378 48832 12384
rect 48410 12271 48466 12280
rect 48228 12096 48280 12102
rect 48228 12038 48280 12044
rect 48320 11892 48372 11898
rect 48320 11834 48372 11840
rect 48332 11150 48360 11834
rect 48320 11144 48372 11150
rect 48320 11086 48372 11092
rect 48228 11008 48280 11014
rect 48226 10976 48228 10985
rect 48280 10976 48282 10985
rect 48226 10911 48282 10920
rect 48136 10056 48188 10062
rect 48136 9998 48188 10004
rect 48148 9450 48176 9998
rect 48136 9444 48188 9450
rect 48136 9386 48188 9392
rect 47584 8832 47636 8838
rect 47584 8774 47636 8780
rect 47768 8832 47820 8838
rect 47768 8774 47820 8780
rect 48136 8832 48188 8838
rect 48136 8774 48188 8780
rect 47596 8498 47624 8774
rect 47584 8492 47636 8498
rect 47584 8434 47636 8440
rect 47596 7954 47624 8434
rect 47584 7948 47636 7954
rect 47584 7890 47636 7896
rect 47596 7410 47624 7890
rect 47676 7880 47728 7886
rect 47674 7848 47676 7857
rect 47728 7848 47730 7857
rect 47674 7783 47730 7792
rect 47584 7404 47636 7410
rect 47584 7346 47636 7352
rect 47584 6792 47636 6798
rect 47584 6734 47636 6740
rect 47676 6792 47728 6798
rect 47676 6734 47728 6740
rect 47596 6390 47624 6734
rect 47584 6384 47636 6390
rect 47688 6361 47716 6734
rect 47584 6326 47636 6332
rect 47674 6352 47730 6361
rect 47674 6287 47730 6296
rect 47780 5710 47808 8774
rect 48148 8498 48176 8774
rect 48136 8492 48188 8498
rect 48136 8434 48188 8440
rect 48136 8288 48188 8294
rect 48136 8230 48188 8236
rect 47860 8084 47912 8090
rect 47860 8026 47912 8032
rect 47872 7886 47900 8026
rect 48148 7886 48176 8230
rect 47860 7880 47912 7886
rect 47860 7822 47912 7828
rect 48136 7880 48188 7886
rect 48136 7822 48188 7828
rect 48148 7546 48176 7822
rect 48240 7818 48268 10911
rect 48320 9512 48372 9518
rect 48320 9454 48372 9460
rect 48332 8838 48360 9454
rect 48320 8832 48372 8838
rect 48320 8774 48372 8780
rect 48320 8628 48372 8634
rect 48320 8570 48372 8576
rect 48332 8537 48360 8570
rect 48318 8528 48374 8537
rect 48318 8463 48374 8472
rect 48320 8424 48372 8430
rect 48320 8366 48372 8372
rect 48332 8265 48360 8366
rect 48318 8256 48374 8265
rect 48318 8191 48374 8200
rect 48424 8090 48452 12271
rect 48516 11898 48544 12310
rect 48700 12294 48820 12322
rect 48596 12232 48648 12238
rect 48594 12200 48596 12209
rect 48648 12200 48650 12209
rect 48594 12135 48650 12144
rect 48596 12096 48648 12102
rect 48596 12038 48648 12044
rect 48504 11892 48556 11898
rect 48504 11834 48556 11840
rect 48608 11762 48636 12038
rect 48596 11756 48648 11762
rect 48596 11698 48648 11704
rect 48688 11756 48740 11762
rect 48688 11698 48740 11704
rect 48504 11552 48556 11558
rect 48504 11494 48556 11500
rect 48516 11150 48544 11494
rect 48504 11144 48556 11150
rect 48504 11086 48556 11092
rect 48516 9489 48544 11086
rect 48608 10033 48636 11698
rect 48700 11354 48728 11698
rect 48792 11694 48820 12294
rect 48780 11688 48832 11694
rect 48780 11630 48832 11636
rect 48780 11552 48832 11558
rect 48780 11494 48832 11500
rect 48688 11348 48740 11354
rect 48688 11290 48740 11296
rect 48792 11150 48820 11494
rect 48780 11144 48832 11150
rect 48780 11086 48832 11092
rect 48884 10674 48912 13824
rect 49068 13802 49096 14214
rect 49056 13796 49108 13802
rect 49056 13738 49108 13744
rect 48964 13728 49016 13734
rect 48964 13670 49016 13676
rect 48976 13462 49004 13670
rect 48964 13456 49016 13462
rect 48964 13398 49016 13404
rect 49054 12608 49110 12617
rect 49054 12543 49110 12552
rect 48962 12336 49018 12345
rect 48962 12271 48964 12280
rect 49016 12271 49018 12280
rect 48964 12242 49016 12248
rect 48964 12164 49016 12170
rect 48964 12106 49016 12112
rect 48976 11830 49004 12106
rect 48964 11824 49016 11830
rect 48964 11766 49016 11772
rect 49068 11354 49096 12543
rect 49160 11898 49188 19178
rect 49712 18834 49740 22510
rect 49804 20534 49832 23054
rect 49792 20528 49844 20534
rect 49792 20470 49844 20476
rect 49700 18828 49752 18834
rect 49700 18770 49752 18776
rect 49516 18148 49568 18154
rect 49516 18090 49568 18096
rect 49528 17678 49556 18090
rect 49792 18080 49844 18086
rect 49792 18022 49844 18028
rect 49804 17746 49832 18022
rect 49792 17740 49844 17746
rect 49792 17682 49844 17688
rect 49516 17672 49568 17678
rect 49516 17614 49568 17620
rect 49332 17264 49384 17270
rect 49332 17206 49384 17212
rect 49238 16416 49294 16425
rect 49238 16351 49294 16360
rect 49252 16250 49280 16351
rect 49240 16244 49292 16250
rect 49240 16186 49292 16192
rect 49238 15464 49294 15473
rect 49238 15399 49240 15408
rect 49292 15399 49294 15408
rect 49240 15370 49292 15376
rect 49344 15026 49372 17206
rect 49424 15972 49476 15978
rect 49424 15914 49476 15920
rect 49332 15020 49384 15026
rect 49332 14962 49384 14968
rect 49330 14920 49386 14929
rect 49330 14855 49332 14864
rect 49384 14855 49386 14864
rect 49332 14826 49384 14832
rect 49332 14408 49384 14414
rect 49332 14350 49384 14356
rect 49344 13841 49372 14350
rect 49436 13870 49464 15914
rect 49528 15473 49556 17614
rect 49608 16516 49660 16522
rect 49608 16458 49660 16464
rect 49514 15464 49570 15473
rect 49514 15399 49570 15408
rect 49516 15360 49568 15366
rect 49516 15302 49568 15308
rect 49424 13864 49476 13870
rect 49330 13832 49386 13841
rect 49424 13806 49476 13812
rect 49330 13767 49386 13776
rect 49240 12806 49292 12812
rect 49240 12748 49292 12754
rect 49148 11892 49200 11898
rect 49148 11834 49200 11840
rect 49148 11688 49200 11694
rect 49148 11630 49200 11636
rect 49056 11348 49108 11354
rect 49056 11290 49108 11296
rect 48872 10668 48924 10674
rect 48872 10610 48924 10616
rect 48884 10198 48912 10610
rect 48872 10192 48924 10198
rect 48778 10160 48834 10169
rect 48688 10124 48740 10130
rect 48872 10134 48924 10140
rect 48778 10095 48834 10104
rect 48688 10066 48740 10072
rect 48594 10024 48650 10033
rect 48594 9959 48650 9968
rect 48596 9716 48648 9722
rect 48596 9658 48648 9664
rect 48502 9480 48558 9489
rect 48502 9415 48558 9424
rect 48516 8974 48544 9415
rect 48504 8968 48556 8974
rect 48504 8910 48556 8916
rect 48412 8084 48464 8090
rect 48412 8026 48464 8032
rect 48228 7812 48280 7818
rect 48228 7754 48280 7760
rect 48136 7540 48188 7546
rect 48136 7482 48188 7488
rect 47860 7268 47912 7274
rect 47860 7210 47912 7216
rect 47768 5704 47820 5710
rect 47768 5646 47820 5652
rect 47492 5636 47544 5642
rect 47492 5578 47544 5584
rect 47136 5528 47256 5556
rect 46940 5510 46992 5516
rect 46664 5364 46716 5370
rect 46848 5364 46900 5370
rect 46716 5324 46796 5352
rect 46664 5306 46716 5312
rect 46570 5264 46626 5273
rect 46570 5199 46626 5208
rect 46480 5024 46532 5030
rect 46480 4966 46532 4972
rect 46662 4720 46718 4729
rect 46662 4655 46718 4664
rect 46676 4554 46704 4655
rect 46664 4548 46716 4554
rect 46664 4490 46716 4496
rect 46388 4480 46440 4486
rect 46388 4422 46440 4428
rect 46204 4276 46256 4282
rect 46204 4218 46256 4224
rect 45928 3392 45980 3398
rect 45928 3334 45980 3340
rect 46216 2650 46244 4218
rect 46480 3936 46532 3942
rect 46480 3878 46532 3884
rect 46492 3602 46520 3878
rect 46480 3596 46532 3602
rect 46480 3538 46532 3544
rect 46664 3460 46716 3466
rect 46664 3402 46716 3408
rect 46676 3126 46704 3402
rect 46768 3126 46796 5324
rect 46848 5306 46900 5312
rect 46952 4622 46980 5510
rect 47032 5228 47084 5234
rect 47032 5170 47084 5176
rect 47044 5001 47072 5170
rect 47030 4992 47086 5001
rect 47030 4927 47086 4936
rect 46940 4616 46992 4622
rect 46940 4558 46992 4564
rect 46664 3120 46716 3126
rect 46664 3062 46716 3068
rect 46756 3120 46808 3126
rect 46756 3062 46808 3068
rect 47228 3058 47256 5528
rect 47504 5370 47532 5578
rect 47492 5364 47544 5370
rect 47492 5306 47544 5312
rect 47872 5302 47900 7210
rect 48240 7002 48268 7754
rect 48412 7472 48464 7478
rect 48412 7414 48464 7420
rect 48228 6996 48280 7002
rect 48228 6938 48280 6944
rect 48318 6896 48374 6905
rect 48318 6831 48374 6840
rect 48044 6792 48096 6798
rect 48044 6734 48096 6740
rect 48056 6322 48084 6734
rect 48044 6316 48096 6322
rect 48044 6258 48096 6264
rect 48056 5710 48084 6258
rect 48332 5846 48360 6831
rect 48320 5840 48372 5846
rect 48320 5782 48372 5788
rect 48044 5704 48096 5710
rect 48044 5646 48096 5652
rect 47860 5296 47912 5302
rect 47860 5238 47912 5244
rect 47674 4992 47730 5001
rect 47674 4927 47730 4936
rect 47398 4856 47454 4865
rect 47688 4826 47716 4927
rect 47398 4791 47400 4800
rect 47452 4791 47454 4800
rect 47676 4820 47728 4826
rect 47400 4762 47452 4768
rect 47676 4762 47728 4768
rect 47768 4752 47820 4758
rect 47768 4694 47820 4700
rect 47308 4480 47360 4486
rect 47492 4480 47544 4486
rect 47360 4440 47492 4468
rect 47308 4422 47360 4428
rect 47492 4422 47544 4428
rect 47582 4448 47638 4457
rect 47582 4383 47638 4392
rect 47596 4214 47624 4383
rect 47584 4208 47636 4214
rect 47584 4150 47636 4156
rect 47596 3738 47624 4150
rect 47584 3732 47636 3738
rect 47584 3674 47636 3680
rect 47780 3194 47808 4694
rect 47872 3670 47900 5238
rect 48044 4548 48096 4554
rect 47964 4508 48044 4536
rect 47964 4457 47992 4508
rect 48044 4490 48096 4496
rect 47950 4448 48006 4457
rect 47950 4383 48006 4392
rect 48136 4004 48188 4010
rect 48136 3946 48188 3952
rect 47860 3664 47912 3670
rect 47860 3606 47912 3612
rect 47768 3188 47820 3194
rect 47768 3130 47820 3136
rect 48148 3126 48176 3946
rect 48228 3936 48280 3942
rect 48228 3878 48280 3884
rect 48136 3120 48188 3126
rect 48136 3062 48188 3068
rect 48240 3058 48268 3878
rect 48424 3126 48452 7414
rect 48608 7410 48636 9658
rect 48700 9654 48728 10066
rect 48688 9648 48740 9654
rect 48688 9590 48740 9596
rect 48792 9568 48820 10095
rect 49056 10056 49108 10062
rect 49056 9998 49108 10004
rect 48872 9580 48924 9586
rect 48792 9540 48872 9568
rect 48686 9344 48742 9353
rect 48686 9279 48742 9288
rect 48596 7404 48648 7410
rect 48596 7346 48648 7352
rect 48596 6996 48648 7002
rect 48596 6938 48648 6944
rect 48608 6322 48636 6938
rect 48700 6730 48728 9279
rect 48688 6724 48740 6730
rect 48688 6666 48740 6672
rect 48596 6316 48648 6322
rect 48596 6258 48648 6264
rect 48608 5710 48636 6258
rect 48792 5914 48820 9540
rect 48872 9522 48924 9528
rect 48964 9444 49016 9450
rect 48964 9386 49016 9392
rect 48976 9217 49004 9386
rect 48962 9208 49018 9217
rect 48962 9143 49018 9152
rect 48872 7404 48924 7410
rect 48872 7346 48924 7352
rect 48964 7404 49016 7410
rect 48964 7346 49016 7352
rect 48884 7041 48912 7346
rect 48870 7032 48926 7041
rect 48870 6967 48926 6976
rect 48780 5908 48832 5914
rect 48780 5850 48832 5856
rect 48780 5772 48832 5778
rect 48780 5714 48832 5720
rect 48596 5704 48648 5710
rect 48596 5646 48648 5652
rect 48608 5234 48636 5646
rect 48688 5636 48740 5642
rect 48688 5578 48740 5584
rect 48596 5228 48648 5234
rect 48596 5170 48648 5176
rect 48502 5128 48558 5137
rect 48502 5063 48504 5072
rect 48556 5063 48558 5072
rect 48504 5034 48556 5040
rect 48596 5024 48648 5030
rect 48596 4966 48648 4972
rect 48608 4486 48636 4966
rect 48596 4480 48648 4486
rect 48596 4422 48648 4428
rect 48412 3120 48464 3126
rect 48412 3062 48464 3068
rect 47216 3052 47268 3058
rect 47216 2994 47268 3000
rect 48228 3052 48280 3058
rect 48228 2994 48280 3000
rect 47124 2984 47176 2990
rect 47124 2926 47176 2932
rect 47030 2680 47086 2689
rect 46204 2644 46256 2650
rect 47030 2615 47032 2624
rect 46204 2586 46256 2592
rect 47084 2615 47086 2624
rect 47032 2586 47084 2592
rect 45652 2576 45704 2582
rect 45652 2518 45704 2524
rect 47044 2446 47072 2586
rect 47136 2582 47164 2926
rect 48700 2650 48728 5578
rect 48792 5030 48820 5714
rect 48780 5024 48832 5030
rect 48780 4966 48832 4972
rect 48792 3126 48820 4966
rect 48872 4684 48924 4690
rect 48872 4626 48924 4632
rect 48884 3534 48912 4626
rect 48976 4214 49004 7346
rect 49068 6866 49096 9998
rect 49160 8838 49188 11630
rect 49252 10266 49280 12748
rect 49240 10260 49292 10266
rect 49240 10202 49292 10208
rect 49344 9722 49372 13767
rect 49422 12880 49478 12889
rect 49422 12815 49424 12824
rect 49476 12815 49478 12824
rect 49424 12786 49476 12792
rect 49424 12368 49476 12374
rect 49528 12356 49556 15302
rect 49620 13734 49648 16458
rect 49700 15972 49752 15978
rect 49700 15914 49752 15920
rect 49608 13728 49660 13734
rect 49606 13696 49608 13705
rect 49660 13696 49662 13705
rect 49606 13631 49662 13640
rect 49712 13433 49740 15914
rect 49792 15156 49844 15162
rect 49792 15098 49844 15104
rect 49804 14550 49832 15098
rect 49792 14544 49844 14550
rect 49792 14486 49844 14492
rect 49698 13424 49754 13433
rect 49698 13359 49700 13368
rect 49752 13359 49754 13368
rect 49700 13330 49752 13336
rect 49792 13320 49844 13326
rect 49792 13262 49844 13268
rect 49700 13252 49752 13258
rect 49700 13194 49752 13200
rect 49608 13184 49660 13190
rect 49608 13126 49660 13132
rect 49620 12986 49648 13126
rect 49608 12980 49660 12986
rect 49608 12922 49660 12928
rect 49608 12640 49660 12646
rect 49608 12582 49660 12588
rect 49476 12328 49556 12356
rect 49424 12310 49476 12316
rect 49620 12238 49648 12582
rect 49712 12306 49740 13194
rect 49804 12918 49832 13262
rect 49896 12986 49924 23718
rect 49976 23724 50028 23730
rect 49976 23666 50028 23672
rect 49988 23254 50016 23666
rect 50172 23322 50200 24550
rect 50724 24410 50752 25298
rect 51000 25294 51028 25842
rect 52196 25838 52224 26206
rect 52184 25832 52236 25838
rect 52184 25774 52236 25780
rect 52380 25362 52408 26930
rect 53208 26858 53236 27814
rect 53760 27470 53788 28018
rect 53748 27464 53800 27470
rect 53748 27406 53800 27412
rect 53196 26852 53248 26858
rect 53196 26794 53248 26800
rect 53380 26784 53432 26790
rect 53380 26726 53432 26732
rect 53392 26586 53420 26726
rect 53380 26580 53432 26586
rect 53380 26522 53432 26528
rect 53852 26382 53880 28358
rect 53944 28014 53972 28562
rect 53932 28008 53984 28014
rect 53932 27950 53984 27956
rect 53944 27470 53972 27950
rect 54128 27470 54156 29106
rect 54208 28076 54260 28082
rect 54208 28018 54260 28024
rect 54392 28076 54444 28082
rect 54392 28018 54444 28024
rect 54220 27606 54248 28018
rect 54208 27600 54260 27606
rect 54208 27542 54260 27548
rect 53932 27464 53984 27470
rect 53932 27406 53984 27412
rect 54116 27464 54168 27470
rect 54116 27406 54168 27412
rect 53944 27334 53972 27406
rect 53932 27328 53984 27334
rect 53932 27270 53984 27276
rect 53840 26376 53892 26382
rect 53840 26318 53892 26324
rect 54024 26376 54076 26382
rect 54024 26318 54076 26324
rect 54036 26042 54064 26318
rect 54024 26036 54076 26042
rect 54024 25978 54076 25984
rect 53196 25900 53248 25906
rect 53196 25842 53248 25848
rect 52736 25832 52788 25838
rect 52736 25774 52788 25780
rect 52460 25696 52512 25702
rect 52460 25638 52512 25644
rect 52368 25356 52420 25362
rect 52368 25298 52420 25304
rect 50988 25288 51040 25294
rect 50988 25230 51040 25236
rect 51000 24954 51028 25230
rect 50988 24948 51040 24954
rect 50988 24890 51040 24896
rect 52472 24818 52500 25638
rect 52748 24886 52776 25774
rect 52828 25356 52880 25362
rect 52828 25298 52880 25304
rect 52736 24880 52788 24886
rect 52736 24822 52788 24828
rect 52460 24812 52512 24818
rect 52460 24754 52512 24760
rect 50712 24404 50764 24410
rect 50712 24346 50764 24352
rect 51632 24268 51684 24274
rect 51632 24210 51684 24216
rect 50804 24200 50856 24206
rect 50804 24142 50856 24148
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50816 23866 50844 24142
rect 50804 23860 50856 23866
rect 50804 23802 50856 23808
rect 51644 23730 51672 24210
rect 52000 23792 52052 23798
rect 52000 23734 52052 23740
rect 51632 23724 51684 23730
rect 51632 23666 51684 23672
rect 50160 23316 50212 23322
rect 50160 23258 50212 23264
rect 49976 23248 50028 23254
rect 49976 23190 50028 23196
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 51264 22636 51316 22642
rect 51264 22578 51316 22584
rect 50160 22092 50212 22098
rect 50160 22034 50212 22040
rect 50068 22024 50120 22030
rect 50068 21966 50120 21972
rect 50080 21690 50108 21966
rect 50068 21684 50120 21690
rect 50068 21626 50120 21632
rect 50080 20466 50108 21626
rect 50172 20466 50200 22034
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 51276 21010 51304 22578
rect 51264 21004 51316 21010
rect 51264 20946 51316 20952
rect 50896 20936 50948 20942
rect 50896 20878 50948 20884
rect 51356 20936 51408 20942
rect 51356 20878 51408 20884
rect 51540 20936 51592 20942
rect 51540 20878 51592 20884
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50908 20534 50936 20878
rect 50896 20528 50948 20534
rect 50896 20470 50948 20476
rect 51080 20528 51132 20534
rect 51080 20470 51132 20476
rect 50068 20460 50120 20466
rect 50068 20402 50120 20408
rect 50160 20460 50212 20466
rect 50160 20402 50212 20408
rect 50172 19514 50200 20402
rect 50908 20398 50936 20470
rect 50896 20392 50948 20398
rect 50896 20334 50948 20340
rect 50908 19854 50936 20334
rect 51092 19854 51120 20470
rect 51172 20460 51224 20466
rect 51172 20402 51224 20408
rect 51184 20058 51212 20402
rect 51172 20052 51224 20058
rect 51172 19994 51224 20000
rect 50896 19848 50948 19854
rect 50896 19790 50948 19796
rect 51080 19848 51132 19854
rect 51080 19790 51132 19796
rect 51080 19712 51132 19718
rect 51080 19654 51132 19660
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50160 19508 50212 19514
rect 50160 19450 50212 19456
rect 50160 19372 50212 19378
rect 50160 19314 50212 19320
rect 49976 19304 50028 19310
rect 49976 19246 50028 19252
rect 49988 16250 50016 19246
rect 50172 18766 50200 19314
rect 50712 19168 50764 19174
rect 50712 19110 50764 19116
rect 50724 18766 50752 19110
rect 51092 18970 51120 19654
rect 51368 19514 51396 20878
rect 51552 20534 51580 20878
rect 51540 20528 51592 20534
rect 51540 20470 51592 20476
rect 51356 19508 51408 19514
rect 51356 19450 51408 19456
rect 51080 18964 51132 18970
rect 51080 18906 51132 18912
rect 50988 18828 51040 18834
rect 50988 18770 51040 18776
rect 50160 18760 50212 18766
rect 50160 18702 50212 18708
rect 50712 18760 50764 18766
rect 50712 18702 50764 18708
rect 50160 18624 50212 18630
rect 50160 18566 50212 18572
rect 50172 18290 50200 18566
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50712 18352 50764 18358
rect 50712 18294 50764 18300
rect 50160 18284 50212 18290
rect 50160 18226 50212 18232
rect 50172 18154 50200 18226
rect 50160 18148 50212 18154
rect 50080 18108 50160 18136
rect 50080 17134 50108 18108
rect 50160 18090 50212 18096
rect 50724 17678 50752 18294
rect 50896 18148 50948 18154
rect 50896 18090 50948 18096
rect 50528 17672 50580 17678
rect 50712 17672 50764 17678
rect 50580 17632 50660 17660
rect 50528 17614 50580 17620
rect 50160 17604 50212 17610
rect 50160 17546 50212 17552
rect 50068 17128 50120 17134
rect 50068 17070 50120 17076
rect 50172 16998 50200 17546
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50434 17232 50490 17241
rect 50434 17167 50436 17176
rect 50488 17167 50490 17176
rect 50436 17138 50488 17144
rect 50526 17096 50582 17105
rect 50526 17031 50582 17040
rect 50160 16992 50212 16998
rect 50160 16934 50212 16940
rect 50068 16584 50120 16590
rect 50068 16526 50120 16532
rect 49976 16244 50028 16250
rect 49976 16186 50028 16192
rect 49976 16040 50028 16046
rect 49976 15982 50028 15988
rect 49988 15609 50016 15982
rect 50080 15638 50108 16526
rect 50172 16232 50200 16934
rect 50540 16590 50568 17031
rect 50528 16584 50580 16590
rect 50528 16526 50580 16532
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50632 16232 50660 17632
rect 50712 17614 50764 17620
rect 50724 17270 50752 17614
rect 50908 17610 50936 18090
rect 51000 17882 51028 18770
rect 51172 18216 51224 18222
rect 51172 18158 51224 18164
rect 51448 18216 51500 18222
rect 51448 18158 51500 18164
rect 50988 17876 51040 17882
rect 50988 17818 51040 17824
rect 50896 17604 50948 17610
rect 50896 17546 50948 17552
rect 50712 17264 50764 17270
rect 50712 17206 50764 17212
rect 50804 16992 50856 16998
rect 50804 16934 50856 16940
rect 50816 16726 50844 16934
rect 50804 16720 50856 16726
rect 50804 16662 50856 16668
rect 50804 16584 50856 16590
rect 50804 16526 50856 16532
rect 50986 16552 51042 16561
rect 50816 16250 50844 16526
rect 50986 16487 51042 16496
rect 51000 16454 51028 16487
rect 50988 16448 51040 16454
rect 50988 16390 51040 16396
rect 50172 16204 50292 16232
rect 50160 16108 50212 16114
rect 50160 16050 50212 16056
rect 50172 15881 50200 16050
rect 50264 15910 50292 16204
rect 50448 16204 50660 16232
rect 50804 16244 50856 16250
rect 50448 16114 50476 16204
rect 50804 16186 50856 16192
rect 50988 16244 51040 16250
rect 50988 16186 51040 16192
rect 50436 16108 50488 16114
rect 50436 16050 50488 16056
rect 50620 16108 50672 16114
rect 50620 16050 50672 16056
rect 50804 16108 50856 16114
rect 50804 16050 50856 16056
rect 50252 15904 50304 15910
rect 50158 15872 50214 15881
rect 50252 15846 50304 15852
rect 50158 15807 50214 15816
rect 50632 15706 50660 16050
rect 50160 15700 50212 15706
rect 50160 15642 50212 15648
rect 50620 15700 50672 15706
rect 50620 15642 50672 15648
rect 50068 15632 50120 15638
rect 49974 15600 50030 15609
rect 50068 15574 50120 15580
rect 49974 15535 50030 15544
rect 49976 15428 50028 15434
rect 49976 15370 50028 15376
rect 49988 15162 50016 15370
rect 49976 15156 50028 15162
rect 49976 15098 50028 15104
rect 49988 14482 50016 15098
rect 50066 15056 50122 15065
rect 50066 14991 50122 15000
rect 50172 15008 50200 15642
rect 50712 15496 50764 15502
rect 50712 15438 50764 15444
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50252 15020 50304 15026
rect 50080 14958 50108 14991
rect 50172 14980 50252 15008
rect 50252 14962 50304 14968
rect 50344 15020 50396 15026
rect 50344 14962 50396 14968
rect 50068 14952 50120 14958
rect 50264 14929 50292 14962
rect 50068 14894 50120 14900
rect 50250 14920 50306 14929
rect 50250 14855 50306 14864
rect 50160 14544 50212 14550
rect 50160 14486 50212 14492
rect 49976 14476 50028 14482
rect 49976 14418 50028 14424
rect 50172 14006 50200 14486
rect 50356 14278 50384 14962
rect 50620 14816 50672 14822
rect 50620 14758 50672 14764
rect 50632 14618 50660 14758
rect 50620 14612 50672 14618
rect 50620 14554 50672 14560
rect 50344 14272 50396 14278
rect 50344 14214 50396 14220
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50160 14000 50212 14006
rect 50160 13942 50212 13948
rect 50172 13870 50200 13942
rect 50620 13932 50672 13938
rect 50620 13874 50672 13880
rect 49976 13864 50028 13870
rect 49976 13806 50028 13812
rect 50160 13864 50212 13870
rect 50160 13806 50212 13812
rect 50436 13864 50488 13870
rect 50436 13806 50488 13812
rect 49884 12980 49936 12986
rect 49884 12922 49936 12928
rect 49792 12912 49844 12918
rect 49844 12860 49924 12866
rect 49792 12854 49924 12860
rect 49804 12838 49924 12854
rect 49792 12776 49844 12782
rect 49792 12718 49844 12724
rect 49700 12300 49752 12306
rect 49700 12242 49752 12248
rect 49608 12232 49660 12238
rect 49608 12174 49660 12180
rect 49424 12096 49476 12102
rect 49424 12038 49476 12044
rect 49436 11558 49464 12038
rect 49516 11688 49568 11694
rect 49516 11630 49568 11636
rect 49424 11552 49476 11558
rect 49424 11494 49476 11500
rect 49528 10538 49556 11630
rect 49698 11112 49754 11121
rect 49698 11047 49700 11056
rect 49752 11047 49754 11056
rect 49700 11018 49752 11024
rect 49700 10600 49752 10606
rect 49700 10542 49752 10548
rect 49516 10532 49568 10538
rect 49516 10474 49568 10480
rect 49424 10464 49476 10470
rect 49424 10406 49476 10412
rect 49514 10432 49570 10441
rect 49436 10266 49464 10406
rect 49514 10367 49570 10376
rect 49424 10260 49476 10266
rect 49424 10202 49476 10208
rect 49424 10056 49476 10062
rect 49422 10024 49424 10033
rect 49476 10024 49478 10033
rect 49422 9959 49478 9968
rect 49332 9716 49384 9722
rect 49332 9658 49384 9664
rect 49240 9648 49292 9654
rect 49240 9590 49292 9596
rect 49252 8974 49280 9590
rect 49240 8968 49292 8974
rect 49240 8910 49292 8916
rect 49148 8832 49200 8838
rect 49148 8774 49200 8780
rect 49056 6860 49108 6866
rect 49056 6802 49108 6808
rect 49160 6390 49188 8774
rect 49528 7886 49556 10367
rect 49608 9104 49660 9110
rect 49608 9046 49660 9052
rect 49620 8906 49648 9046
rect 49608 8900 49660 8906
rect 49608 8842 49660 8848
rect 49606 8528 49662 8537
rect 49606 8463 49608 8472
rect 49660 8463 49662 8472
rect 49608 8434 49660 8440
rect 49712 8378 49740 10542
rect 49804 10470 49832 12718
rect 49792 10464 49844 10470
rect 49790 10432 49792 10441
rect 49844 10432 49846 10441
rect 49790 10367 49846 10376
rect 49792 9988 49844 9994
rect 49792 9930 49844 9936
rect 49804 9586 49832 9930
rect 49792 9580 49844 9586
rect 49792 9522 49844 9528
rect 49792 9104 49844 9110
rect 49792 9046 49844 9052
rect 49804 8634 49832 9046
rect 49792 8628 49844 8634
rect 49792 8570 49844 8576
rect 49620 8350 49740 8378
rect 49792 8424 49844 8430
rect 49792 8366 49844 8372
rect 49332 7880 49384 7886
rect 49332 7822 49384 7828
rect 49516 7880 49568 7886
rect 49516 7822 49568 7828
rect 49344 7721 49372 7822
rect 49330 7712 49386 7721
rect 49330 7647 49386 7656
rect 49620 7449 49648 8350
rect 49700 8288 49752 8294
rect 49700 8230 49752 8236
rect 49606 7440 49662 7449
rect 49606 7375 49662 7384
rect 49620 7342 49648 7375
rect 49608 7336 49660 7342
rect 49608 7278 49660 7284
rect 49332 7268 49384 7274
rect 49332 7210 49384 7216
rect 49344 6798 49372 7210
rect 49424 7200 49476 7206
rect 49424 7142 49476 7148
rect 49436 7002 49464 7142
rect 49424 6996 49476 7002
rect 49424 6938 49476 6944
rect 49332 6792 49384 6798
rect 49332 6734 49384 6740
rect 49712 6746 49740 8230
rect 49804 7954 49832 8366
rect 49896 8090 49924 12838
rect 49988 12714 50016 13806
rect 50448 13530 50476 13806
rect 50068 13524 50120 13530
rect 50068 13466 50120 13472
rect 50436 13524 50488 13530
rect 50436 13466 50488 13472
rect 49976 12708 50028 12714
rect 49976 12650 50028 12656
rect 49976 12232 50028 12238
rect 49976 12174 50028 12180
rect 49988 11150 50016 12174
rect 49976 11144 50028 11150
rect 49976 11086 50028 11092
rect 50080 11082 50108 13466
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50632 12968 50660 13874
rect 50724 13326 50752 15438
rect 50712 13320 50764 13326
rect 50712 13262 50764 13268
rect 50448 12940 50660 12968
rect 50342 12608 50398 12617
rect 50342 12543 50398 12552
rect 50356 12306 50384 12543
rect 50344 12300 50396 12306
rect 50344 12242 50396 12248
rect 50448 12170 50476 12940
rect 50620 12844 50672 12850
rect 50620 12786 50672 12792
rect 50436 12164 50488 12170
rect 50436 12106 50488 12112
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50632 11898 50660 12786
rect 50712 12436 50764 12442
rect 50712 12378 50764 12384
rect 50620 11892 50672 11898
rect 50620 11834 50672 11840
rect 50724 11286 50752 12378
rect 50816 12209 50844 16050
rect 50896 15020 50948 15026
rect 50896 14962 50948 14968
rect 50908 14521 50936 14962
rect 50894 14512 50950 14521
rect 50894 14447 50950 14456
rect 51000 13682 51028 16186
rect 51184 16182 51212 18158
rect 51356 17536 51408 17542
rect 51356 17478 51408 17484
rect 51368 17202 51396 17478
rect 51460 17338 51488 18158
rect 51448 17332 51500 17338
rect 51448 17274 51500 17280
rect 51356 17196 51408 17202
rect 51264 17158 51316 17164
rect 51356 17138 51408 17144
rect 51264 17100 51316 17106
rect 51172 16176 51224 16182
rect 51276 16153 51304 17100
rect 51356 16584 51408 16590
rect 51354 16552 51356 16561
rect 51408 16552 51410 16561
rect 51354 16487 51410 16496
rect 51540 16516 51592 16522
rect 51540 16458 51592 16464
rect 51552 16250 51580 16458
rect 51540 16244 51592 16250
rect 51540 16186 51592 16192
rect 51172 16118 51224 16124
rect 51262 16144 51318 16153
rect 51080 15972 51132 15978
rect 51080 15914 51132 15920
rect 51092 14822 51120 15914
rect 51080 14816 51132 14822
rect 51080 14758 51132 14764
rect 51184 14618 51212 16118
rect 51262 16079 51318 16088
rect 51540 16108 51592 16114
rect 51276 15094 51304 16079
rect 51540 16050 51592 16056
rect 51356 16040 51408 16046
rect 51356 15982 51408 15988
rect 51264 15088 51316 15094
rect 51264 15030 51316 15036
rect 51172 14612 51224 14618
rect 51172 14554 51224 14560
rect 51172 14408 51224 14414
rect 51172 14350 51224 14356
rect 51184 13802 51212 14350
rect 51264 13932 51316 13938
rect 51264 13874 51316 13880
rect 51172 13796 51224 13802
rect 51172 13738 51224 13744
rect 50908 13654 51028 13682
rect 50802 12200 50858 12209
rect 50802 12135 50858 12144
rect 50804 12096 50856 12102
rect 50804 12038 50856 12044
rect 50816 11898 50844 12038
rect 50804 11892 50856 11898
rect 50804 11834 50856 11840
rect 50908 11354 50936 13654
rect 50988 13524 51040 13530
rect 50988 13466 51040 13472
rect 51000 12782 51028 13466
rect 51172 13184 51224 13190
rect 51172 13126 51224 13132
rect 50988 12776 51040 12782
rect 50988 12718 51040 12724
rect 51080 12708 51132 12714
rect 51080 12650 51132 12656
rect 50986 12064 51042 12073
rect 50986 11999 51042 12008
rect 50896 11348 50948 11354
rect 50896 11290 50948 11296
rect 50712 11280 50764 11286
rect 50764 11240 50844 11268
rect 50712 11222 50764 11228
rect 50160 11144 50212 11150
rect 50160 11086 50212 11092
rect 50528 11144 50580 11150
rect 50528 11086 50580 11092
rect 50816 11098 50844 11240
rect 51000 11234 51028 11999
rect 51092 11830 51120 12650
rect 51080 11824 51132 11830
rect 51080 11766 51132 11772
rect 51080 11280 51132 11286
rect 51000 11228 51080 11234
rect 51000 11222 51132 11228
rect 51000 11206 51120 11222
rect 51080 11144 51132 11150
rect 50068 11076 50120 11082
rect 50068 11018 50120 11024
rect 50172 10674 50200 11086
rect 50540 11014 50568 11086
rect 50816 11070 51028 11098
rect 51080 11086 51132 11092
rect 50528 11008 50580 11014
rect 50528 10950 50580 10956
rect 50712 11008 50764 11014
rect 50712 10950 50764 10956
rect 50896 11008 50948 11014
rect 50896 10950 50948 10956
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50160 10668 50212 10674
rect 50160 10610 50212 10616
rect 50172 10198 50200 10610
rect 50528 10600 50580 10606
rect 50528 10542 50580 10548
rect 50540 10282 50568 10542
rect 50436 10260 50488 10266
rect 50540 10254 50660 10282
rect 50436 10202 50488 10208
rect 50160 10192 50212 10198
rect 50160 10134 50212 10140
rect 50068 9580 50120 9586
rect 50068 9522 50120 9528
rect 49976 9376 50028 9382
rect 49976 9318 50028 9324
rect 49988 8974 50016 9318
rect 50080 9217 50108 9522
rect 50066 9208 50122 9217
rect 50066 9143 50122 9152
rect 50068 9036 50120 9042
rect 50068 8978 50120 8984
rect 49976 8968 50028 8974
rect 49976 8910 50028 8916
rect 49884 8084 49936 8090
rect 49884 8026 49936 8032
rect 49792 7948 49844 7954
rect 49792 7890 49844 7896
rect 49884 7812 49936 7818
rect 49884 7754 49936 7760
rect 49792 7744 49844 7750
rect 49896 7721 49924 7754
rect 49792 7686 49844 7692
rect 49882 7712 49938 7721
rect 49804 7410 49832 7686
rect 49882 7647 49938 7656
rect 49792 7404 49844 7410
rect 49792 7346 49844 7352
rect 49896 7342 49924 7647
rect 49884 7336 49936 7342
rect 49884 7278 49936 7284
rect 49792 7200 49844 7206
rect 49792 7142 49844 7148
rect 49804 6866 49832 7142
rect 49792 6860 49844 6866
rect 49792 6802 49844 6808
rect 49884 6792 49936 6798
rect 49790 6760 49846 6769
rect 49712 6718 49790 6746
rect 49884 6734 49936 6740
rect 49790 6695 49846 6704
rect 49148 6384 49200 6390
rect 49148 6326 49200 6332
rect 49804 6118 49832 6695
rect 49896 6458 49924 6734
rect 49884 6452 49936 6458
rect 49884 6394 49936 6400
rect 49884 6248 49936 6254
rect 49884 6190 49936 6196
rect 49792 6112 49844 6118
rect 49792 6054 49844 6060
rect 49606 5808 49662 5817
rect 49896 5778 49924 6190
rect 49606 5743 49662 5752
rect 49884 5772 49936 5778
rect 49620 5710 49648 5743
rect 49884 5714 49936 5720
rect 49608 5704 49660 5710
rect 49608 5646 49660 5652
rect 49698 5672 49754 5681
rect 49332 5228 49384 5234
rect 49332 5170 49384 5176
rect 49056 5160 49108 5166
rect 49240 5160 49292 5166
rect 49108 5120 49240 5148
rect 49056 5102 49108 5108
rect 49240 5102 49292 5108
rect 49344 4690 49372 5170
rect 49620 5166 49648 5646
rect 49698 5607 49754 5616
rect 49712 5370 49740 5607
rect 49700 5364 49752 5370
rect 49700 5306 49752 5312
rect 49608 5160 49660 5166
rect 49608 5102 49660 5108
rect 49332 4684 49384 4690
rect 49332 4626 49384 4632
rect 49608 4480 49660 4486
rect 49608 4422 49660 4428
rect 49620 4214 49648 4422
rect 48964 4208 49016 4214
rect 48964 4150 49016 4156
rect 49608 4208 49660 4214
rect 49608 4150 49660 4156
rect 49896 4146 49924 5714
rect 49988 4758 50016 8910
rect 50080 8498 50108 8978
rect 50068 8492 50120 8498
rect 50068 8434 50120 8440
rect 50172 8430 50200 10134
rect 50448 10062 50476 10202
rect 50436 10056 50488 10062
rect 50436 9998 50488 10004
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50252 9648 50304 9654
rect 50252 9590 50304 9596
rect 50264 9178 50292 9590
rect 50252 9172 50304 9178
rect 50252 9114 50304 9120
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50252 8560 50304 8566
rect 50632 8537 50660 10254
rect 50724 9926 50752 10950
rect 50908 10198 50936 10950
rect 50896 10192 50948 10198
rect 50896 10134 50948 10140
rect 50804 10056 50856 10062
rect 50804 9998 50856 10004
rect 50712 9920 50764 9926
rect 50712 9862 50764 9868
rect 50724 8634 50752 9862
rect 50816 9178 50844 9998
rect 51000 9674 51028 11070
rect 51092 10810 51120 11086
rect 51080 10804 51132 10810
rect 51080 10746 51132 10752
rect 50908 9654 51028 9674
rect 50896 9648 51028 9654
rect 50948 9646 51028 9648
rect 50896 9590 50948 9596
rect 50908 9438 51120 9466
rect 50804 9172 50856 9178
rect 50804 9114 50856 9120
rect 50908 8838 50936 9438
rect 51092 9382 51120 9438
rect 51080 9376 51132 9382
rect 51080 9318 51132 9324
rect 51184 8838 51212 13126
rect 51276 12345 51304 13874
rect 51368 13530 51396 15982
rect 51448 15904 51500 15910
rect 51552 15881 51580 16050
rect 51448 15846 51500 15852
rect 51538 15872 51594 15881
rect 51460 15162 51488 15846
rect 51538 15807 51594 15816
rect 51644 15706 51672 23666
rect 51908 23520 51960 23526
rect 51908 23462 51960 23468
rect 51724 22636 51776 22642
rect 51724 22578 51776 22584
rect 51736 17882 51764 22578
rect 51816 20256 51868 20262
rect 51816 20198 51868 20204
rect 51724 17876 51776 17882
rect 51724 17818 51776 17824
rect 51828 17678 51856 20198
rect 51920 18902 51948 23462
rect 52012 22982 52040 23734
rect 52092 23724 52144 23730
rect 52092 23666 52144 23672
rect 52184 23724 52236 23730
rect 52184 23666 52236 23672
rect 52104 23322 52132 23666
rect 52092 23316 52144 23322
rect 52092 23258 52144 23264
rect 52000 22976 52052 22982
rect 52000 22918 52052 22924
rect 52012 22778 52040 22918
rect 52000 22772 52052 22778
rect 52000 22714 52052 22720
rect 52104 22574 52132 23258
rect 52196 23118 52224 23666
rect 52472 23526 52500 24754
rect 52748 24206 52776 24822
rect 52840 24800 52868 25298
rect 53208 24818 53236 25842
rect 54220 25770 54248 27542
rect 54404 27538 54432 28018
rect 55232 28014 55260 29106
rect 57152 28552 57204 28558
rect 57152 28494 57204 28500
rect 56968 28416 57020 28422
rect 56968 28358 57020 28364
rect 55588 28076 55640 28082
rect 55588 28018 55640 28024
rect 55864 28076 55916 28082
rect 55864 28018 55916 28024
rect 56048 28076 56100 28082
rect 56048 28018 56100 28024
rect 55220 28008 55272 28014
rect 55220 27950 55272 27956
rect 54392 27532 54444 27538
rect 54392 27474 54444 27480
rect 54404 27130 54432 27474
rect 55232 27470 55260 27950
rect 55600 27606 55628 28018
rect 55588 27600 55640 27606
rect 55588 27542 55640 27548
rect 54576 27464 54628 27470
rect 54576 27406 54628 27412
rect 55220 27464 55272 27470
rect 55220 27406 55272 27412
rect 54392 27124 54444 27130
rect 54392 27066 54444 27072
rect 54588 27062 54616 27406
rect 54576 27056 54628 27062
rect 54576 26998 54628 27004
rect 55876 26994 55904 28018
rect 56060 26994 56088 28018
rect 56980 27470 57008 28358
rect 56968 27464 57020 27470
rect 56968 27406 57020 27412
rect 57164 27130 57192 28494
rect 57244 28484 57296 28490
rect 57244 28426 57296 28432
rect 57256 28150 57284 28426
rect 57244 28144 57296 28150
rect 57244 28086 57296 28092
rect 57152 27124 57204 27130
rect 57152 27066 57204 27072
rect 54300 26988 54352 26994
rect 54300 26930 54352 26936
rect 54944 26988 54996 26994
rect 55864 26988 55916 26994
rect 54944 26930 54996 26936
rect 55784 26948 55864 26976
rect 54312 25906 54340 26930
rect 54956 26518 54984 26930
rect 55220 26784 55272 26790
rect 55220 26726 55272 26732
rect 54944 26512 54996 26518
rect 54944 26454 54996 26460
rect 54300 25900 54352 25906
rect 54300 25842 54352 25848
rect 54392 25900 54444 25906
rect 54392 25842 54444 25848
rect 54208 25764 54260 25770
rect 54208 25706 54260 25712
rect 53288 25696 53340 25702
rect 53288 25638 53340 25644
rect 53300 25294 53328 25638
rect 54312 25498 54340 25842
rect 54300 25492 54352 25498
rect 54300 25434 54352 25440
rect 54404 25362 54432 25842
rect 54392 25356 54444 25362
rect 54392 25298 54444 25304
rect 53288 25288 53340 25294
rect 53288 25230 53340 25236
rect 53932 25288 53984 25294
rect 53932 25230 53984 25236
rect 54208 25288 54260 25294
rect 54208 25230 54260 25236
rect 53944 24818 53972 25230
rect 52920 24812 52972 24818
rect 52840 24772 52920 24800
rect 52920 24754 52972 24760
rect 53196 24812 53248 24818
rect 53196 24754 53248 24760
rect 53932 24812 53984 24818
rect 53932 24754 53984 24760
rect 52736 24200 52788 24206
rect 52736 24142 52788 24148
rect 52552 24132 52604 24138
rect 52552 24074 52604 24080
rect 52460 23520 52512 23526
rect 52460 23462 52512 23468
rect 52184 23112 52236 23118
rect 52184 23054 52236 23060
rect 52196 22574 52224 23054
rect 52092 22568 52144 22574
rect 52092 22510 52144 22516
rect 52184 22568 52236 22574
rect 52184 22510 52236 22516
rect 52564 21078 52592 24074
rect 52644 22500 52696 22506
rect 52644 22442 52696 22448
rect 52656 21962 52684 22442
rect 52644 21956 52696 21962
rect 52644 21898 52696 21904
rect 52828 21956 52880 21962
rect 52828 21898 52880 21904
rect 52840 21690 52868 21898
rect 52828 21684 52880 21690
rect 52828 21626 52880 21632
rect 52552 21072 52604 21078
rect 52552 21014 52604 21020
rect 52000 21004 52052 21010
rect 52000 20946 52052 20952
rect 52012 19854 52040 20946
rect 52564 20466 52592 21014
rect 52552 20460 52604 20466
rect 52552 20402 52604 20408
rect 52736 20392 52788 20398
rect 52736 20334 52788 20340
rect 52748 19854 52776 20334
rect 52828 19916 52880 19922
rect 52828 19858 52880 19864
rect 52000 19848 52052 19854
rect 52000 19790 52052 19796
rect 52736 19848 52788 19854
rect 52736 19790 52788 19796
rect 52012 19446 52040 19790
rect 52092 19712 52144 19718
rect 52092 19654 52144 19660
rect 52104 19514 52132 19654
rect 52092 19508 52144 19514
rect 52092 19450 52144 19456
rect 52000 19440 52052 19446
rect 52000 19382 52052 19388
rect 52000 19304 52052 19310
rect 51998 19272 52000 19281
rect 52052 19272 52054 19281
rect 51998 19207 52054 19216
rect 51908 18896 51960 18902
rect 51908 18838 51960 18844
rect 52460 18760 52512 18766
rect 52460 18702 52512 18708
rect 52184 18420 52236 18426
rect 52184 18362 52236 18368
rect 51908 18284 51960 18290
rect 51908 18226 51960 18232
rect 51920 18086 51948 18226
rect 51908 18080 51960 18086
rect 51908 18022 51960 18028
rect 51816 17672 51868 17678
rect 51816 17614 51868 17620
rect 51920 17542 51948 18022
rect 52196 17746 52224 18362
rect 52368 18080 52420 18086
rect 52368 18022 52420 18028
rect 52184 17740 52236 17746
rect 52184 17682 52236 17688
rect 52000 17672 52052 17678
rect 52000 17614 52052 17620
rect 51908 17536 51960 17542
rect 51908 17478 51960 17484
rect 51920 17134 51948 17478
rect 52012 17202 52040 17614
rect 52000 17196 52052 17202
rect 52000 17138 52052 17144
rect 51908 17128 51960 17134
rect 51908 17070 51960 17076
rect 51632 15700 51684 15706
rect 51632 15642 51684 15648
rect 51816 15632 51868 15638
rect 51816 15574 51868 15580
rect 51448 15156 51500 15162
rect 51448 15098 51500 15104
rect 51448 15020 51500 15026
rect 51448 14962 51500 14968
rect 51724 15020 51776 15026
rect 51724 14962 51776 14968
rect 51356 13524 51408 13530
rect 51356 13466 51408 13472
rect 51356 13388 51408 13394
rect 51356 13330 51408 13336
rect 51368 12782 51396 13330
rect 51460 13190 51488 14962
rect 51632 14952 51684 14958
rect 51632 14894 51684 14900
rect 51540 14340 51592 14346
rect 51540 14282 51592 14288
rect 51552 14006 51580 14282
rect 51540 14000 51592 14006
rect 51540 13942 51592 13948
rect 51644 13938 51672 14894
rect 51632 13932 51684 13938
rect 51632 13874 51684 13880
rect 51448 13184 51500 13190
rect 51448 13126 51500 13132
rect 51356 12776 51408 12782
rect 51356 12718 51408 12724
rect 51368 12434 51396 12718
rect 51368 12406 51488 12434
rect 51262 12336 51318 12345
rect 51262 12271 51318 12280
rect 51356 11620 51408 11626
rect 51356 11562 51408 11568
rect 51368 10606 51396 11562
rect 51356 10600 51408 10606
rect 51356 10542 51408 10548
rect 51356 10464 51408 10470
rect 51356 10406 51408 10412
rect 51368 10062 51396 10406
rect 51460 10198 51488 12406
rect 51644 12356 51672 13874
rect 51736 12434 51764 14962
rect 51828 13394 51856 15574
rect 51920 15570 51948 17070
rect 52012 16998 52040 17138
rect 52000 16992 52052 16998
rect 52000 16934 52052 16940
rect 52000 16108 52052 16114
rect 52000 16050 52052 16056
rect 51908 15564 51960 15570
rect 51908 15506 51960 15512
rect 51906 14784 51962 14793
rect 51906 14719 51962 14728
rect 51920 14618 51948 14719
rect 51908 14612 51960 14618
rect 51908 14554 51960 14560
rect 51920 14414 51948 14554
rect 51908 14408 51960 14414
rect 51908 14350 51960 14356
rect 52012 13444 52040 16050
rect 52196 14618 52224 17682
rect 52380 17678 52408 18022
rect 52368 17672 52420 17678
rect 52368 17614 52420 17620
rect 52368 17128 52420 17134
rect 52368 17070 52420 17076
rect 52276 16788 52328 16794
rect 52276 16730 52328 16736
rect 52288 16522 52316 16730
rect 52276 16516 52328 16522
rect 52276 16458 52328 16464
rect 52276 15496 52328 15502
rect 52276 15438 52328 15444
rect 52380 15484 52408 17070
rect 52472 15858 52500 18702
rect 52840 18426 52868 19858
rect 52932 18834 52960 24754
rect 53012 24336 53064 24342
rect 53012 24278 53064 24284
rect 53024 23730 53052 24278
rect 53104 24200 53156 24206
rect 53104 24142 53156 24148
rect 53116 23866 53144 24142
rect 53104 23860 53156 23866
rect 53104 23802 53156 23808
rect 53012 23724 53064 23730
rect 53012 23666 53064 23672
rect 53024 23050 53052 23666
rect 53208 23322 53236 24754
rect 53932 24200 53984 24206
rect 53932 24142 53984 24148
rect 53288 23724 53340 23730
rect 53288 23666 53340 23672
rect 53840 23724 53892 23730
rect 53840 23666 53892 23672
rect 53300 23322 53328 23666
rect 53852 23322 53880 23666
rect 53944 23662 53972 24142
rect 54220 23866 54248 25230
rect 54760 24812 54812 24818
rect 54760 24754 54812 24760
rect 54668 24200 54720 24206
rect 54668 24142 54720 24148
rect 54208 23860 54260 23866
rect 54208 23802 54260 23808
rect 53932 23656 53984 23662
rect 53932 23598 53984 23604
rect 53196 23316 53248 23322
rect 53196 23258 53248 23264
rect 53288 23316 53340 23322
rect 53288 23258 53340 23264
rect 53840 23316 53892 23322
rect 53840 23258 53892 23264
rect 53012 23044 53064 23050
rect 53012 22986 53064 22992
rect 53196 23044 53248 23050
rect 53196 22986 53248 22992
rect 53104 22228 53156 22234
rect 53104 22170 53156 22176
rect 53116 21962 53144 22170
rect 53104 21956 53156 21962
rect 53104 21898 53156 21904
rect 53012 20936 53064 20942
rect 53012 20878 53064 20884
rect 53024 20262 53052 20878
rect 53208 20398 53236 22986
rect 53300 22234 53328 23258
rect 53380 22636 53432 22642
rect 53380 22578 53432 22584
rect 53564 22636 53616 22642
rect 53564 22578 53616 22584
rect 53748 22636 53800 22642
rect 53748 22578 53800 22584
rect 53288 22228 53340 22234
rect 53288 22170 53340 22176
rect 53392 22030 53420 22578
rect 53576 22098 53604 22578
rect 53656 22568 53708 22574
rect 53656 22510 53708 22516
rect 53564 22092 53616 22098
rect 53564 22034 53616 22040
rect 53668 22030 53696 22510
rect 53760 22030 53788 22578
rect 53380 22024 53432 22030
rect 53380 21966 53432 21972
rect 53656 22024 53708 22030
rect 53656 21966 53708 21972
rect 53748 22024 53800 22030
rect 53748 21966 53800 21972
rect 53668 21842 53696 21966
rect 53668 21814 53880 21842
rect 53852 20942 53880 21814
rect 53288 20936 53340 20942
rect 53288 20878 53340 20884
rect 53840 20936 53892 20942
rect 53840 20878 53892 20884
rect 53300 20602 53328 20878
rect 53288 20596 53340 20602
rect 53288 20538 53340 20544
rect 53196 20392 53248 20398
rect 53196 20334 53248 20340
rect 53012 20256 53064 20262
rect 53012 20198 53064 20204
rect 52920 18828 52972 18834
rect 52920 18770 52972 18776
rect 52828 18420 52880 18426
rect 52828 18362 52880 18368
rect 52828 17808 52880 17814
rect 52828 17750 52880 17756
rect 52736 17740 52788 17746
rect 52736 17682 52788 17688
rect 52748 17270 52776 17682
rect 52840 17270 52868 17750
rect 53024 17338 53052 20198
rect 53564 19916 53616 19922
rect 53564 19858 53616 19864
rect 53104 19848 53156 19854
rect 53104 19790 53156 19796
rect 53116 19514 53144 19790
rect 53288 19780 53340 19786
rect 53288 19722 53340 19728
rect 53104 19508 53156 19514
rect 53104 19450 53156 19456
rect 53300 19174 53328 19722
rect 53380 19712 53432 19718
rect 53380 19654 53432 19660
rect 53392 19378 53420 19654
rect 53380 19372 53432 19378
rect 53380 19314 53432 19320
rect 53576 19310 53604 19858
rect 53564 19304 53616 19310
rect 53564 19246 53616 19252
rect 53288 19168 53340 19174
rect 53288 19110 53340 19116
rect 53656 19168 53708 19174
rect 53656 19110 53708 19116
rect 53104 17876 53156 17882
rect 53104 17818 53156 17824
rect 53012 17332 53064 17338
rect 53012 17274 53064 17280
rect 52736 17264 52788 17270
rect 52736 17206 52788 17212
rect 52828 17264 52880 17270
rect 53116 17241 53144 17818
rect 53196 17672 53248 17678
rect 53196 17614 53248 17620
rect 52828 17206 52880 17212
rect 53102 17232 53158 17241
rect 52748 16998 52776 17206
rect 53012 17196 53064 17202
rect 53102 17167 53158 17176
rect 53012 17138 53064 17144
rect 52736 16992 52788 16998
rect 52736 16934 52788 16940
rect 52552 16652 52604 16658
rect 52552 16594 52604 16600
rect 52564 16454 52592 16594
rect 52644 16584 52696 16590
rect 52644 16526 52696 16532
rect 52552 16448 52604 16454
rect 52552 16390 52604 16396
rect 52564 16017 52592 16390
rect 52550 16008 52606 16017
rect 52550 15943 52606 15952
rect 52472 15830 52592 15858
rect 52460 15496 52512 15502
rect 52380 15456 52460 15484
rect 52288 14890 52316 15438
rect 52276 14884 52328 14890
rect 52276 14826 52328 14832
rect 52184 14612 52236 14618
rect 52184 14554 52236 14560
rect 52380 14498 52408 15456
rect 52460 15438 52512 15444
rect 52458 15056 52514 15065
rect 52458 14991 52514 15000
rect 52288 14470 52408 14498
rect 52472 14498 52500 14991
rect 52564 14618 52592 15830
rect 52552 14612 52604 14618
rect 52552 14554 52604 14560
rect 52472 14470 52592 14498
rect 52656 14482 52684 16526
rect 52288 14414 52316 14470
rect 52092 14408 52144 14414
rect 52092 14350 52144 14356
rect 52276 14408 52328 14414
rect 52276 14350 52328 14356
rect 52104 14074 52132 14350
rect 52276 14272 52328 14278
rect 52276 14214 52328 14220
rect 52092 14068 52144 14074
rect 52092 14010 52144 14016
rect 52288 13938 52316 14214
rect 52380 14074 52408 14470
rect 52460 14408 52512 14414
rect 52460 14350 52512 14356
rect 52368 14068 52420 14074
rect 52368 14010 52420 14016
rect 52472 13954 52500 14350
rect 52276 13932 52328 13938
rect 52276 13874 52328 13880
rect 52380 13926 52500 13954
rect 52184 13796 52236 13802
rect 52184 13738 52236 13744
rect 52196 13530 52224 13738
rect 52184 13524 52236 13530
rect 52184 13466 52236 13472
rect 52012 13416 52132 13444
rect 51816 13388 51868 13394
rect 51868 13348 52040 13376
rect 51816 13330 51868 13336
rect 51908 12844 51960 12850
rect 51908 12786 51960 12792
rect 51736 12406 51856 12434
rect 51644 12328 51764 12356
rect 51632 12164 51684 12170
rect 51632 12106 51684 12112
rect 51644 11694 51672 12106
rect 51632 11688 51684 11694
rect 51632 11630 51684 11636
rect 51736 11558 51764 12328
rect 51724 11552 51776 11558
rect 51724 11494 51776 11500
rect 51540 11144 51592 11150
rect 51540 11086 51592 11092
rect 51552 10198 51580 11086
rect 51632 11076 51684 11082
rect 51632 11018 51684 11024
rect 51644 10674 51672 11018
rect 51724 10736 51776 10742
rect 51724 10678 51776 10684
rect 51632 10668 51684 10674
rect 51632 10610 51684 10616
rect 51644 10266 51672 10610
rect 51632 10260 51684 10266
rect 51632 10202 51684 10208
rect 51736 10198 51764 10678
rect 51448 10192 51500 10198
rect 51448 10134 51500 10140
rect 51540 10192 51592 10198
rect 51540 10134 51592 10140
rect 51724 10192 51776 10198
rect 51724 10134 51776 10140
rect 51356 10056 51408 10062
rect 51356 9998 51408 10004
rect 51356 9104 51408 9110
rect 51356 9046 51408 9052
rect 50896 8832 50948 8838
rect 50896 8774 50948 8780
rect 51172 8832 51224 8838
rect 51172 8774 51224 8780
rect 50712 8628 50764 8634
rect 50712 8570 50764 8576
rect 50252 8502 50304 8508
rect 50618 8528 50674 8537
rect 50160 8424 50212 8430
rect 50160 8366 50212 8372
rect 50068 7948 50120 7954
rect 50068 7890 50120 7896
rect 50080 7546 50108 7890
rect 50264 7732 50292 8502
rect 50908 8514 50936 8774
rect 50618 8463 50674 8472
rect 50724 8486 50936 8514
rect 50620 8356 50672 8362
rect 50620 8298 50672 8304
rect 50172 7704 50292 7732
rect 50068 7540 50120 7546
rect 50068 7482 50120 7488
rect 50080 6186 50108 7482
rect 50172 6934 50200 7704
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50160 6928 50212 6934
rect 50160 6870 50212 6876
rect 50172 6322 50200 6870
rect 50344 6792 50396 6798
rect 50342 6760 50344 6769
rect 50396 6760 50398 6769
rect 50342 6695 50398 6704
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50344 6452 50396 6458
rect 50344 6394 50396 6400
rect 50356 6361 50384 6394
rect 50342 6352 50398 6361
rect 50160 6316 50212 6322
rect 50342 6287 50344 6296
rect 50160 6258 50212 6264
rect 50396 6287 50398 6296
rect 50344 6258 50396 6264
rect 50436 6248 50488 6254
rect 50436 6190 50488 6196
rect 50068 6180 50120 6186
rect 50068 6122 50120 6128
rect 49976 4752 50028 4758
rect 49976 4694 50028 4700
rect 49884 4140 49936 4146
rect 49884 4082 49936 4088
rect 50080 3738 50108 6122
rect 50448 5914 50476 6190
rect 50436 5908 50488 5914
rect 50436 5850 50488 5856
rect 50632 5846 50660 8298
rect 50724 6322 50752 8486
rect 50804 8424 50856 8430
rect 50804 8366 50856 8372
rect 50816 8090 50844 8366
rect 50896 8288 50948 8294
rect 50896 8230 50948 8236
rect 50988 8288 51040 8294
rect 50988 8230 51040 8236
rect 50804 8084 50856 8090
rect 50804 8026 50856 8032
rect 50816 7002 50844 8026
rect 50804 6996 50856 7002
rect 50804 6938 50856 6944
rect 50804 6792 50856 6798
rect 50804 6734 50856 6740
rect 50816 6390 50844 6734
rect 50804 6384 50856 6390
rect 50804 6326 50856 6332
rect 50712 6316 50764 6322
rect 50712 6258 50764 6264
rect 50620 5840 50672 5846
rect 50620 5782 50672 5788
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50528 5296 50580 5302
rect 50528 5238 50580 5244
rect 50540 4622 50568 5238
rect 50632 5098 50660 5782
rect 50620 5092 50672 5098
rect 50620 5034 50672 5040
rect 50160 4616 50212 4622
rect 50160 4558 50212 4564
rect 50528 4616 50580 4622
rect 50528 4558 50580 4564
rect 50068 3732 50120 3738
rect 50068 3674 50120 3680
rect 49240 3664 49292 3670
rect 49240 3606 49292 3612
rect 48872 3528 48924 3534
rect 48872 3470 48924 3476
rect 48780 3120 48832 3126
rect 48780 3062 48832 3068
rect 48884 2650 48912 3470
rect 49252 3398 49280 3606
rect 49240 3392 49292 3398
rect 49240 3334 49292 3340
rect 48688 2644 48740 2650
rect 48688 2586 48740 2592
rect 48872 2644 48924 2650
rect 48872 2586 48924 2592
rect 49252 2582 49280 3334
rect 50172 3126 50200 4558
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50724 4010 50752 6258
rect 50816 5370 50844 6326
rect 50908 5710 50936 8230
rect 51000 7954 51028 8230
rect 51184 8022 51212 8774
rect 51368 8634 51396 9046
rect 51356 8628 51408 8634
rect 51356 8570 51408 8576
rect 51460 8566 51488 10134
rect 51552 9489 51580 10134
rect 51632 10056 51684 10062
rect 51632 9998 51684 10004
rect 51538 9480 51594 9489
rect 51538 9415 51594 9424
rect 51552 9110 51580 9415
rect 51540 9104 51592 9110
rect 51540 9046 51592 9052
rect 51448 8560 51500 8566
rect 51354 8528 51410 8537
rect 51448 8502 51500 8508
rect 51354 8463 51410 8472
rect 51368 8412 51396 8463
rect 51448 8424 51500 8430
rect 51368 8384 51448 8412
rect 51448 8366 51500 8372
rect 51540 8424 51592 8430
rect 51540 8366 51592 8372
rect 51172 8016 51224 8022
rect 51172 7958 51224 7964
rect 51356 8016 51408 8022
rect 51356 7958 51408 7964
rect 50988 7948 51040 7954
rect 50988 7890 51040 7896
rect 51080 7744 51132 7750
rect 51080 7686 51132 7692
rect 51092 7342 51120 7686
rect 51184 7562 51212 7958
rect 51184 7534 51304 7562
rect 51276 7478 51304 7534
rect 51264 7472 51316 7478
rect 51264 7414 51316 7420
rect 51368 7410 51396 7958
rect 51460 7818 51488 8366
rect 51552 7886 51580 8366
rect 51540 7880 51592 7886
rect 51540 7822 51592 7828
rect 51448 7812 51500 7818
rect 51448 7754 51500 7760
rect 51356 7404 51408 7410
rect 51356 7346 51408 7352
rect 51080 7336 51132 7342
rect 51078 7304 51080 7313
rect 51132 7304 51134 7313
rect 51368 7290 51396 7346
rect 51078 7239 51134 7248
rect 51276 7262 51396 7290
rect 51092 6848 51120 7239
rect 51276 6934 51304 7262
rect 51264 6928 51316 6934
rect 51264 6870 51316 6876
rect 51000 6820 51120 6848
rect 51000 5914 51028 6820
rect 51460 6390 51488 7754
rect 51552 7546 51580 7822
rect 51644 7750 51672 9998
rect 51724 8900 51776 8906
rect 51724 8842 51776 8848
rect 51632 7744 51684 7750
rect 51632 7686 51684 7692
rect 51540 7540 51592 7546
rect 51540 7482 51592 7488
rect 51736 7206 51764 8842
rect 51828 8276 51856 12406
rect 51920 9654 51948 12786
rect 52012 11898 52040 13348
rect 52104 12918 52132 13416
rect 52092 12912 52144 12918
rect 52092 12854 52144 12860
rect 52104 12714 52132 12854
rect 52092 12708 52144 12714
rect 52092 12650 52144 12656
rect 52104 12442 52132 12650
rect 52092 12436 52144 12442
rect 52092 12378 52144 12384
rect 52184 12232 52236 12238
rect 52184 12174 52236 12180
rect 52000 11892 52052 11898
rect 52000 11834 52052 11840
rect 52092 11620 52144 11626
rect 52092 11562 52144 11568
rect 52000 11144 52052 11150
rect 52000 11086 52052 11092
rect 52012 10810 52040 11086
rect 52104 11082 52132 11562
rect 52196 11354 52224 12174
rect 52184 11348 52236 11354
rect 52184 11290 52236 11296
rect 52182 11248 52238 11257
rect 52182 11183 52238 11192
rect 52092 11076 52144 11082
rect 52092 11018 52144 11024
rect 52000 10804 52052 10810
rect 52000 10746 52052 10752
rect 52196 10674 52224 11183
rect 52092 10668 52144 10674
rect 52092 10610 52144 10616
rect 52184 10668 52236 10674
rect 52184 10610 52236 10616
rect 52000 10192 52052 10198
rect 52000 10134 52052 10140
rect 51908 9648 51960 9654
rect 51908 9590 51960 9596
rect 52012 9058 52040 10134
rect 52104 9722 52132 10610
rect 52196 10577 52224 10610
rect 52182 10568 52238 10577
rect 52182 10503 52238 10512
rect 52184 10260 52236 10266
rect 52184 10202 52236 10208
rect 52092 9716 52144 9722
rect 52092 9658 52144 9664
rect 51920 9030 52040 9058
rect 51920 8430 51948 9030
rect 51908 8424 51960 8430
rect 51908 8366 51960 8372
rect 51828 8248 51948 8276
rect 51814 8120 51870 8129
rect 51814 8055 51816 8064
rect 51868 8055 51870 8064
rect 51816 8026 51868 8032
rect 51920 7954 51948 8248
rect 52104 8090 52132 9658
rect 52196 9625 52224 10202
rect 52182 9616 52238 9625
rect 52182 9551 52238 9560
rect 52184 8492 52236 8498
rect 52184 8434 52236 8440
rect 52092 8084 52144 8090
rect 52092 8026 52144 8032
rect 51908 7948 51960 7954
rect 51908 7890 51960 7896
rect 52000 7880 52052 7886
rect 52196 7868 52224 8434
rect 52288 8022 52316 13874
rect 52380 13569 52408 13926
rect 52366 13560 52422 13569
rect 52366 13495 52422 13504
rect 52564 13512 52592 14470
rect 52644 14476 52696 14482
rect 52644 14418 52696 14424
rect 52748 14414 52776 16934
rect 53024 16726 53052 17138
rect 53012 16720 53064 16726
rect 53012 16662 53064 16668
rect 53116 16658 53144 17167
rect 53208 16697 53236 17614
rect 53194 16688 53250 16697
rect 53104 16652 53156 16658
rect 53194 16623 53250 16632
rect 53104 16594 53156 16600
rect 53196 16516 53248 16522
rect 53196 16458 53248 16464
rect 53208 15502 53236 16458
rect 53196 15496 53248 15502
rect 53196 15438 53248 15444
rect 52920 15428 52972 15434
rect 52920 15370 52972 15376
rect 52828 15360 52880 15366
rect 52828 15302 52880 15308
rect 52840 15094 52868 15302
rect 52828 15088 52880 15094
rect 52828 15030 52880 15036
rect 52932 14618 52960 15370
rect 53012 15088 53064 15094
rect 53012 15030 53064 15036
rect 52920 14612 52972 14618
rect 52920 14554 52972 14560
rect 53024 14532 53052 15030
rect 53104 14544 53156 14550
rect 53024 14504 53104 14532
rect 52736 14408 52788 14414
rect 52736 14350 52788 14356
rect 52828 13864 52880 13870
rect 52828 13806 52880 13812
rect 52840 13530 52868 13806
rect 52920 13728 52972 13734
rect 52920 13670 52972 13676
rect 52828 13524 52880 13530
rect 52380 12730 52408 13495
rect 52564 13484 52776 13512
rect 52644 13388 52696 13394
rect 52644 13330 52696 13336
rect 52460 13320 52512 13326
rect 52460 13262 52512 13268
rect 52472 12850 52500 13262
rect 52552 13184 52604 13190
rect 52552 13126 52604 13132
rect 52564 12918 52592 13126
rect 52552 12912 52604 12918
rect 52552 12854 52604 12860
rect 52460 12844 52512 12850
rect 52460 12786 52512 12792
rect 52380 12702 52500 12730
rect 52368 12232 52420 12238
rect 52366 12200 52368 12209
rect 52420 12200 52422 12209
rect 52366 12135 52422 12144
rect 52368 11756 52420 11762
rect 52368 11698 52420 11704
rect 52380 10985 52408 11698
rect 52366 10976 52422 10985
rect 52366 10911 52422 10920
rect 52472 10826 52500 12702
rect 52564 12238 52592 12854
rect 52552 12232 52604 12238
rect 52552 12174 52604 12180
rect 52552 11892 52604 11898
rect 52552 11834 52604 11840
rect 52564 11014 52592 11834
rect 52552 11008 52604 11014
rect 52552 10950 52604 10956
rect 52380 10798 52500 10826
rect 52276 8016 52328 8022
rect 52276 7958 52328 7964
rect 52052 7840 52224 7868
rect 52000 7822 52052 7828
rect 51724 7200 51776 7206
rect 51724 7142 51776 7148
rect 51736 6798 51764 7142
rect 51724 6792 51776 6798
rect 51724 6734 51776 6740
rect 51908 6792 51960 6798
rect 51908 6734 51960 6740
rect 51540 6452 51592 6458
rect 51540 6394 51592 6400
rect 51448 6384 51500 6390
rect 51170 6352 51226 6361
rect 51448 6326 51500 6332
rect 51170 6287 51172 6296
rect 51224 6287 51226 6296
rect 51172 6258 51224 6264
rect 51552 6186 51580 6394
rect 51736 6361 51764 6734
rect 51722 6352 51778 6361
rect 51722 6287 51724 6296
rect 51776 6287 51778 6296
rect 51724 6258 51776 6264
rect 51736 6227 51764 6258
rect 51540 6180 51592 6186
rect 51540 6122 51592 6128
rect 50988 5908 51040 5914
rect 50988 5850 51040 5856
rect 51920 5778 51948 6734
rect 51908 5772 51960 5778
rect 51908 5714 51960 5720
rect 50896 5704 50948 5710
rect 50896 5646 50948 5652
rect 50804 5364 50856 5370
rect 50804 5306 50856 5312
rect 50804 5024 50856 5030
rect 50804 4966 50856 4972
rect 50816 4690 50844 4966
rect 50804 4684 50856 4690
rect 50804 4626 50856 4632
rect 50908 4146 50936 5646
rect 51538 5264 51594 5273
rect 51538 5199 51594 5208
rect 51632 5228 51684 5234
rect 51552 4826 51580 5199
rect 51632 5170 51684 5176
rect 51644 5030 51672 5170
rect 51632 5024 51684 5030
rect 51632 4966 51684 4972
rect 51540 4820 51592 4826
rect 51540 4762 51592 4768
rect 51644 4593 51672 4966
rect 51630 4584 51686 4593
rect 52012 4554 52040 7822
rect 52288 7426 52316 7958
rect 52196 7410 52316 7426
rect 52184 7404 52316 7410
rect 52236 7398 52316 7404
rect 52184 7346 52236 7352
rect 52276 6792 52328 6798
rect 52276 6734 52328 6740
rect 52288 6390 52316 6734
rect 52184 6384 52236 6390
rect 52184 6326 52236 6332
rect 52276 6384 52328 6390
rect 52276 6326 52328 6332
rect 52196 6254 52224 6326
rect 52184 6248 52236 6254
rect 52184 6190 52236 6196
rect 51630 4519 51686 4528
rect 52000 4548 52052 4554
rect 50896 4140 50948 4146
rect 50896 4082 50948 4088
rect 50712 4004 50764 4010
rect 50712 3946 50764 3952
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50724 3126 50752 3946
rect 50908 3194 50936 4082
rect 51172 3936 51224 3942
rect 51172 3878 51224 3884
rect 51184 3670 51212 3878
rect 51172 3664 51224 3670
rect 51172 3606 51224 3612
rect 51448 3528 51500 3534
rect 51448 3470 51500 3476
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 50896 3188 50948 3194
rect 50896 3130 50948 3136
rect 50160 3120 50212 3126
rect 50160 3062 50212 3068
rect 50712 3120 50764 3126
rect 50712 3062 50764 3068
rect 50908 2650 50936 3130
rect 51368 3058 51396 3402
rect 51460 3194 51488 3470
rect 51448 3188 51500 3194
rect 51448 3130 51500 3136
rect 51356 3052 51408 3058
rect 51356 2994 51408 3000
rect 51644 2650 51672 4519
rect 52000 4490 52052 4496
rect 52012 3466 52040 4490
rect 52196 4010 52224 6190
rect 52288 5234 52316 6326
rect 52380 5914 52408 10798
rect 52460 10600 52512 10606
rect 52460 10542 52512 10548
rect 52472 9761 52500 10542
rect 52656 10470 52684 13330
rect 52748 12374 52776 13484
rect 52828 13466 52880 13472
rect 52736 12368 52788 12374
rect 52736 12310 52788 12316
rect 52748 11665 52776 12310
rect 52840 12238 52868 13466
rect 52932 12850 52960 13670
rect 52920 12844 52972 12850
rect 52920 12786 52972 12792
rect 53024 12458 53052 14504
rect 53104 14486 53156 14492
rect 53104 14272 53156 14278
rect 53104 14214 53156 14220
rect 53116 13297 53144 14214
rect 53208 13326 53236 15438
rect 53300 15162 53328 19110
rect 53668 18290 53696 19110
rect 53944 18698 53972 23598
rect 54680 23050 54708 24142
rect 54772 24138 54800 24754
rect 54760 24132 54812 24138
rect 54760 24074 54812 24080
rect 54668 23044 54720 23050
rect 54668 22986 54720 22992
rect 54680 22710 54708 22986
rect 54668 22704 54720 22710
rect 54668 22646 54720 22652
rect 54392 21956 54444 21962
rect 54392 21898 54444 21904
rect 54300 21888 54352 21894
rect 54300 21830 54352 21836
rect 54404 21842 54432 21898
rect 54312 20942 54340 21830
rect 54404 21814 54708 21842
rect 54404 21690 54432 21814
rect 54392 21684 54444 21690
rect 54392 21626 54444 21632
rect 54484 21616 54536 21622
rect 54484 21558 54536 21564
rect 54392 21548 54444 21554
rect 54392 21490 54444 21496
rect 54404 21146 54432 21490
rect 54392 21140 54444 21146
rect 54392 21082 54444 21088
rect 54024 20936 54076 20942
rect 54024 20878 54076 20884
rect 54300 20936 54352 20942
rect 54300 20878 54352 20884
rect 54036 20466 54064 20878
rect 54024 20460 54076 20466
rect 54024 20402 54076 20408
rect 54208 20460 54260 20466
rect 54208 20402 54260 20408
rect 54220 20058 54248 20402
rect 54312 20262 54340 20878
rect 54496 20482 54524 21558
rect 54576 21344 54628 21350
rect 54576 21286 54628 21292
rect 54588 20942 54616 21286
rect 54576 20936 54628 20942
rect 54576 20878 54628 20884
rect 54404 20466 54524 20482
rect 54404 20460 54536 20466
rect 54404 20454 54484 20460
rect 54300 20256 54352 20262
rect 54300 20198 54352 20204
rect 54208 20052 54260 20058
rect 54208 19994 54260 20000
rect 54024 19984 54076 19990
rect 54404 19938 54432 20454
rect 54484 20402 54536 20408
rect 54484 20324 54536 20330
rect 54484 20266 54536 20272
rect 54024 19926 54076 19932
rect 54036 19718 54064 19926
rect 54128 19910 54432 19938
rect 54128 19854 54156 19910
rect 54496 19854 54524 20266
rect 54116 19848 54168 19854
rect 54116 19790 54168 19796
rect 54300 19848 54352 19854
rect 54300 19790 54352 19796
rect 54484 19848 54536 19854
rect 54484 19790 54536 19796
rect 54024 19712 54076 19718
rect 54024 19654 54076 19660
rect 54116 19372 54168 19378
rect 54116 19314 54168 19320
rect 54024 18760 54076 18766
rect 54024 18702 54076 18708
rect 53932 18692 53984 18698
rect 53932 18634 53984 18640
rect 53748 18352 53800 18358
rect 53748 18294 53800 18300
rect 53656 18284 53708 18290
rect 53656 18226 53708 18232
rect 53472 17876 53524 17882
rect 53472 17818 53524 17824
rect 53484 16794 53512 17818
rect 53668 17134 53696 18226
rect 53656 17128 53708 17134
rect 53656 17070 53708 17076
rect 53760 16794 53788 18294
rect 53932 18284 53984 18290
rect 53932 18226 53984 18232
rect 53840 17672 53892 17678
rect 53840 17614 53892 17620
rect 53852 17202 53880 17614
rect 53944 17338 53972 18226
rect 54036 18057 54064 18702
rect 54022 18048 54078 18057
rect 54022 17983 54078 17992
rect 54128 17678 54156 19314
rect 54208 18148 54260 18154
rect 54208 18090 54260 18096
rect 54116 17672 54168 17678
rect 54116 17614 54168 17620
rect 53932 17332 53984 17338
rect 53932 17274 53984 17280
rect 54128 17270 54156 17614
rect 54220 17542 54248 18090
rect 54208 17536 54260 17542
rect 54208 17478 54260 17484
rect 54116 17264 54168 17270
rect 54116 17206 54168 17212
rect 53840 17196 53892 17202
rect 53840 17138 53892 17144
rect 53932 17196 53984 17202
rect 53932 17138 53984 17144
rect 53472 16788 53524 16794
rect 53472 16730 53524 16736
rect 53748 16788 53800 16794
rect 53748 16730 53800 16736
rect 53840 16652 53892 16658
rect 53840 16594 53892 16600
rect 53380 16584 53432 16590
rect 53380 16526 53432 16532
rect 53288 15156 53340 15162
rect 53288 15098 53340 15104
rect 53288 14952 53340 14958
rect 53288 14894 53340 14900
rect 53300 14414 53328 14894
rect 53288 14408 53340 14414
rect 53288 14350 53340 14356
rect 53392 14074 53420 16526
rect 53748 16448 53800 16454
rect 53748 16390 53800 16396
rect 53760 16046 53788 16390
rect 53852 16114 53880 16594
rect 53840 16108 53892 16114
rect 53840 16050 53892 16056
rect 53748 16040 53800 16046
rect 53748 15982 53800 15988
rect 53472 15496 53524 15502
rect 53472 15438 53524 15444
rect 53484 14929 53512 15438
rect 53656 15360 53708 15366
rect 53656 15302 53708 15308
rect 53470 14920 53526 14929
rect 53470 14855 53472 14864
rect 53524 14855 53526 14864
rect 53472 14826 53524 14832
rect 53484 14795 53512 14826
rect 53380 14068 53432 14074
rect 53380 14010 53432 14016
rect 53288 13864 53340 13870
rect 53288 13806 53340 13812
rect 53196 13320 53248 13326
rect 53102 13288 53158 13297
rect 53196 13262 53248 13268
rect 53102 13223 53158 13232
rect 53116 12850 53144 13223
rect 53196 13184 53248 13190
rect 53196 13126 53248 13132
rect 53104 12844 53156 12850
rect 53104 12786 53156 12792
rect 53024 12430 53144 12458
rect 52828 12232 52880 12238
rect 52828 12174 52880 12180
rect 52734 11656 52790 11665
rect 52734 11591 52790 11600
rect 52736 11552 52788 11558
rect 52736 11494 52788 11500
rect 52644 10464 52696 10470
rect 52644 10406 52696 10412
rect 52656 10266 52684 10406
rect 52644 10260 52696 10266
rect 52644 10202 52696 10208
rect 52458 9752 52514 9761
rect 52458 9687 52514 9696
rect 52748 9654 52776 11494
rect 52736 9648 52788 9654
rect 52458 9616 52514 9625
rect 52736 9590 52788 9596
rect 52458 9551 52460 9560
rect 52512 9551 52514 9560
rect 52460 9522 52512 9528
rect 52472 6866 52500 9522
rect 52552 9512 52604 9518
rect 52840 9500 52868 12174
rect 52920 12164 52972 12170
rect 52920 12106 52972 12112
rect 52932 10674 52960 12106
rect 53116 11150 53144 12430
rect 53208 12186 53236 13126
rect 53300 12306 53328 13806
rect 53380 13796 53432 13802
rect 53380 13738 53432 13744
rect 53392 12434 53420 13738
rect 53472 13320 53524 13326
rect 53472 13262 53524 13268
rect 53484 12730 53512 13262
rect 53668 13190 53696 15302
rect 53760 13394 53788 15982
rect 53840 15360 53892 15366
rect 53840 15302 53892 15308
rect 53852 15065 53880 15302
rect 53838 15056 53894 15065
rect 53838 14991 53894 15000
rect 53840 14408 53892 14414
rect 53840 14350 53892 14356
rect 53748 13388 53800 13394
rect 53748 13330 53800 13336
rect 53656 13184 53708 13190
rect 53656 13126 53708 13132
rect 53852 12986 53880 14350
rect 53944 13870 53972 17138
rect 54128 16250 54156 17206
rect 54208 17128 54260 17134
rect 54208 17070 54260 17076
rect 54116 16244 54168 16250
rect 54116 16186 54168 16192
rect 54024 15020 54076 15026
rect 54128 15008 54156 16186
rect 54220 16046 54248 17070
rect 54312 16561 54340 19790
rect 54496 17882 54524 19790
rect 54484 17876 54536 17882
rect 54484 17818 54536 17824
rect 54484 17536 54536 17542
rect 54484 17478 54536 17484
rect 54496 17134 54524 17478
rect 54588 17338 54616 20878
rect 54576 17332 54628 17338
rect 54576 17274 54628 17280
rect 54680 17218 54708 21814
rect 54772 20534 54800 24074
rect 54760 20528 54812 20534
rect 54760 20470 54812 20476
rect 54760 20256 54812 20262
rect 54760 20198 54812 20204
rect 54772 19922 54800 20198
rect 54760 19916 54812 19922
rect 54760 19858 54812 19864
rect 54956 19514 54984 26454
rect 55036 25900 55088 25906
rect 55036 25842 55088 25848
rect 55048 25294 55076 25842
rect 55232 25702 55260 26726
rect 55220 25696 55272 25702
rect 55220 25638 55272 25644
rect 55036 25288 55088 25294
rect 55036 25230 55088 25236
rect 55496 24812 55548 24818
rect 55496 24754 55548 24760
rect 55508 24206 55536 24754
rect 55784 24274 55812 26948
rect 56048 26988 56100 26994
rect 55864 26930 55916 26936
rect 55968 26948 56048 26976
rect 55968 26314 55996 26948
rect 56048 26930 56100 26936
rect 56968 26988 57020 26994
rect 56968 26930 57020 26936
rect 56324 26920 56376 26926
rect 56324 26862 56376 26868
rect 56336 26382 56364 26862
rect 56980 26518 57008 26930
rect 57060 26852 57112 26858
rect 57060 26794 57112 26800
rect 56508 26512 56560 26518
rect 56508 26454 56560 26460
rect 56968 26512 57020 26518
rect 56968 26454 57020 26460
rect 56520 26382 56548 26454
rect 56324 26376 56376 26382
rect 56324 26318 56376 26324
rect 56508 26376 56560 26382
rect 56508 26318 56560 26324
rect 55956 26308 56008 26314
rect 55956 26250 56008 26256
rect 56336 26234 56364 26318
rect 57072 26314 57100 26794
rect 57060 26308 57112 26314
rect 57060 26250 57112 26256
rect 56336 26206 56456 26234
rect 56048 25900 56100 25906
rect 56100 25860 56180 25888
rect 56048 25842 56100 25848
rect 55864 25832 55916 25838
rect 55864 25774 55916 25780
rect 55876 25294 55904 25774
rect 55956 25696 56008 25702
rect 55956 25638 56008 25644
rect 55968 25498 55996 25638
rect 55956 25492 56008 25498
rect 55956 25434 56008 25440
rect 56152 25362 56180 25860
rect 56140 25356 56192 25362
rect 56140 25298 56192 25304
rect 55864 25288 55916 25294
rect 55864 25230 55916 25236
rect 55876 24410 55904 25230
rect 55864 24404 55916 24410
rect 55864 24346 55916 24352
rect 55772 24268 55824 24274
rect 55772 24210 55824 24216
rect 55496 24200 55548 24206
rect 55496 24142 55548 24148
rect 55128 22636 55180 22642
rect 55128 22578 55180 22584
rect 55036 21956 55088 21962
rect 55036 21898 55088 21904
rect 55048 21554 55076 21898
rect 55140 21894 55168 22578
rect 55220 22024 55272 22030
rect 55220 21966 55272 21972
rect 55128 21888 55180 21894
rect 55128 21830 55180 21836
rect 55140 21690 55168 21830
rect 55128 21684 55180 21690
rect 55128 21626 55180 21632
rect 55232 21554 55260 21966
rect 55036 21548 55088 21554
rect 55036 21490 55088 21496
rect 55220 21548 55272 21554
rect 55220 21490 55272 21496
rect 55232 20602 55260 21490
rect 55508 21078 55536 24142
rect 56152 23254 56180 25298
rect 56324 24812 56376 24818
rect 56324 24754 56376 24760
rect 56336 24070 56364 24754
rect 56428 24750 56456 26206
rect 57072 25906 57100 26250
rect 57164 26042 57192 27066
rect 57256 26926 57284 28086
rect 57244 26920 57296 26926
rect 57244 26862 57296 26868
rect 57152 26036 57204 26042
rect 57152 25978 57204 25984
rect 57060 25900 57112 25906
rect 57060 25842 57112 25848
rect 57152 25900 57204 25906
rect 57256 25888 57284 26862
rect 57204 25860 57284 25888
rect 57152 25842 57204 25848
rect 56876 25696 56928 25702
rect 56876 25638 56928 25644
rect 56416 24744 56468 24750
rect 56416 24686 56468 24692
rect 56508 24744 56560 24750
rect 56508 24686 56560 24692
rect 56416 24200 56468 24206
rect 56416 24142 56468 24148
rect 56324 24064 56376 24070
rect 56324 24006 56376 24012
rect 56336 23730 56364 24006
rect 56428 23866 56456 24142
rect 56416 23860 56468 23866
rect 56416 23802 56468 23808
rect 56520 23746 56548 24686
rect 56888 24138 56916 25638
rect 57072 25498 57100 25842
rect 57060 25492 57112 25498
rect 57060 25434 57112 25440
rect 57060 25220 57112 25226
rect 57060 25162 57112 25168
rect 56968 24608 57020 24614
rect 56968 24550 57020 24556
rect 56980 24206 57008 24550
rect 56968 24200 57020 24206
rect 56968 24142 57020 24148
rect 56876 24132 56928 24138
rect 56876 24074 56928 24080
rect 56428 23730 56548 23746
rect 56324 23724 56376 23730
rect 56324 23666 56376 23672
rect 56416 23724 56548 23730
rect 56468 23718 56548 23724
rect 56416 23666 56468 23672
rect 56428 23610 56456 23666
rect 56336 23582 56456 23610
rect 56888 23594 56916 24074
rect 56876 23588 56928 23594
rect 56140 23248 56192 23254
rect 56140 23190 56192 23196
rect 55588 23180 55640 23186
rect 55588 23122 55640 23128
rect 55600 22642 55628 23122
rect 55680 23112 55732 23118
rect 55680 23054 55732 23060
rect 55588 22636 55640 22642
rect 55588 22578 55640 22584
rect 55496 21072 55548 21078
rect 55496 21014 55548 21020
rect 55404 21004 55456 21010
rect 55404 20946 55456 20952
rect 55220 20596 55272 20602
rect 55220 20538 55272 20544
rect 55416 20466 55444 20946
rect 55404 20460 55456 20466
rect 55404 20402 55456 20408
rect 55416 19786 55444 20402
rect 55496 19848 55548 19854
rect 55496 19790 55548 19796
rect 55404 19780 55456 19786
rect 55404 19722 55456 19728
rect 55508 19718 55536 19790
rect 55496 19712 55548 19718
rect 55496 19654 55548 19660
rect 54944 19508 54996 19514
rect 54944 19450 54996 19456
rect 55496 19304 55548 19310
rect 55496 19246 55548 19252
rect 55508 18970 55536 19246
rect 55496 18964 55548 18970
rect 55496 18906 55548 18912
rect 55128 18760 55180 18766
rect 55128 18702 55180 18708
rect 55140 18426 55168 18702
rect 55128 18420 55180 18426
rect 55128 18362 55180 18368
rect 54760 18080 54812 18086
rect 54760 18022 54812 18028
rect 54588 17190 54708 17218
rect 54484 17128 54536 17134
rect 54484 17070 54536 17076
rect 54298 16552 54354 16561
rect 54298 16487 54354 16496
rect 54484 16516 54536 16522
rect 54208 16040 54260 16046
rect 54208 15982 54260 15988
rect 54208 15020 54260 15026
rect 54128 14980 54208 15008
rect 54024 14962 54076 14968
rect 54208 14962 54260 14968
rect 53932 13864 53984 13870
rect 53932 13806 53984 13812
rect 53840 12980 53892 12986
rect 53840 12922 53892 12928
rect 53748 12776 53800 12782
rect 53484 12702 53696 12730
rect 53748 12718 53800 12724
rect 53564 12640 53616 12646
rect 53564 12582 53616 12588
rect 53392 12406 53512 12434
rect 53380 12368 53432 12374
rect 53378 12336 53380 12345
rect 53432 12336 53434 12345
rect 53288 12300 53340 12306
rect 53378 12271 53434 12280
rect 53288 12242 53340 12248
rect 53208 12158 53328 12186
rect 53196 11824 53248 11830
rect 53196 11766 53248 11772
rect 53012 11144 53064 11150
rect 53104 11144 53156 11150
rect 53012 11086 53064 11092
rect 53102 11112 53104 11121
rect 53156 11112 53158 11121
rect 53024 10742 53052 11086
rect 53102 11047 53158 11056
rect 53104 11008 53156 11014
rect 53104 10950 53156 10956
rect 53012 10736 53064 10742
rect 53012 10678 53064 10684
rect 52920 10668 52972 10674
rect 52920 10610 52972 10616
rect 53116 10266 53144 10950
rect 53104 10260 53156 10266
rect 53104 10202 53156 10208
rect 53012 10124 53064 10130
rect 53012 10066 53064 10072
rect 52920 9648 52972 9654
rect 52920 9590 52972 9596
rect 52552 9454 52604 9460
rect 52748 9472 52868 9500
rect 52564 9353 52592 9454
rect 52550 9344 52606 9353
rect 52606 9302 52684 9330
rect 52550 9279 52606 9288
rect 52552 9036 52604 9042
rect 52552 8978 52604 8984
rect 52564 8945 52592 8978
rect 52656 8974 52684 9302
rect 52644 8968 52696 8974
rect 52550 8936 52606 8945
rect 52644 8910 52696 8916
rect 52550 8871 52606 8880
rect 52656 7750 52684 8910
rect 52748 8906 52776 9472
rect 52932 8922 52960 9590
rect 53024 9450 53052 10066
rect 53104 10056 53156 10062
rect 53104 9998 53156 10004
rect 53116 9926 53144 9998
rect 53104 9920 53156 9926
rect 53104 9862 53156 9868
rect 53012 9444 53064 9450
rect 53012 9386 53064 9392
rect 53116 8922 53144 9862
rect 52736 8900 52788 8906
rect 52736 8842 52788 8848
rect 52840 8894 53144 8922
rect 53208 9568 53236 11766
rect 53300 11626 53328 12158
rect 53380 11688 53432 11694
rect 53380 11630 53432 11636
rect 53288 11620 53340 11626
rect 53288 11562 53340 11568
rect 53300 11082 53328 11562
rect 53288 11076 53340 11082
rect 53288 11018 53340 11024
rect 53300 10674 53328 11018
rect 53288 10668 53340 10674
rect 53288 10610 53340 10616
rect 53300 10198 53328 10610
rect 53288 10192 53340 10198
rect 53288 10134 53340 10140
rect 53288 9580 53340 9586
rect 53208 9540 53288 9568
rect 52644 7744 52696 7750
rect 52644 7686 52696 7692
rect 52552 7540 52604 7546
rect 52552 7482 52604 7488
rect 52736 7540 52788 7546
rect 52736 7482 52788 7488
rect 52460 6860 52512 6866
rect 52460 6802 52512 6808
rect 52460 6724 52512 6730
rect 52460 6666 52512 6672
rect 52472 6254 52500 6666
rect 52564 6662 52592 7482
rect 52748 7206 52776 7482
rect 52736 7200 52788 7206
rect 52736 7142 52788 7148
rect 52840 6934 52868 8894
rect 53012 8832 53064 8838
rect 53012 8774 53064 8780
rect 53024 8634 53052 8774
rect 53208 8634 53236 9540
rect 53288 9522 53340 9528
rect 53012 8628 53064 8634
rect 53012 8570 53064 8576
rect 53196 8628 53248 8634
rect 53196 8570 53248 8576
rect 52920 8492 52972 8498
rect 52920 8434 52972 8440
rect 52932 7410 52960 8434
rect 53024 7886 53052 8570
rect 53012 7880 53064 7886
rect 53012 7822 53064 7828
rect 53288 7880 53340 7886
rect 53288 7822 53340 7828
rect 52920 7404 52972 7410
rect 52920 7346 52972 7352
rect 52932 7002 52960 7346
rect 52920 6996 52972 7002
rect 52920 6938 52972 6944
rect 52828 6928 52880 6934
rect 52828 6870 52880 6876
rect 52552 6656 52604 6662
rect 52552 6598 52604 6604
rect 52736 6656 52788 6662
rect 52736 6598 52788 6604
rect 52460 6248 52512 6254
rect 52460 6190 52512 6196
rect 52368 5908 52420 5914
rect 52368 5850 52420 5856
rect 52276 5228 52328 5234
rect 52276 5170 52328 5176
rect 52184 4004 52236 4010
rect 52184 3946 52236 3952
rect 52000 3460 52052 3466
rect 52000 3402 52052 3408
rect 51908 3188 51960 3194
rect 51908 3130 51960 3136
rect 51920 2650 51948 3130
rect 52196 3058 52224 3946
rect 52288 3534 52316 5170
rect 52564 4214 52592 6598
rect 52748 6390 52776 6598
rect 52736 6384 52788 6390
rect 52736 6326 52788 6332
rect 52840 4826 52868 6870
rect 53024 6254 53052 7822
rect 53300 7342 53328 7822
rect 53288 7336 53340 7342
rect 53288 7278 53340 7284
rect 53300 6730 53328 7278
rect 53392 7206 53420 11630
rect 53484 9926 53512 12406
rect 53576 12238 53604 12582
rect 53668 12442 53696 12702
rect 53656 12436 53708 12442
rect 53656 12378 53708 12384
rect 53656 12300 53708 12306
rect 53656 12242 53708 12248
rect 53564 12232 53616 12238
rect 53668 12209 53696 12242
rect 53564 12174 53616 12180
rect 53654 12200 53710 12209
rect 53654 12135 53710 12144
rect 53564 12096 53616 12102
rect 53564 12038 53616 12044
rect 53576 11762 53604 12038
rect 53564 11756 53616 11762
rect 53564 11698 53616 11704
rect 53564 11008 53616 11014
rect 53564 10950 53616 10956
rect 53472 9920 53524 9926
rect 53472 9862 53524 9868
rect 53470 9752 53526 9761
rect 53470 9687 53526 9696
rect 53484 9586 53512 9687
rect 53472 9580 53524 9586
rect 53472 9522 53524 9528
rect 53472 7948 53524 7954
rect 53472 7890 53524 7896
rect 53484 7410 53512 7890
rect 53472 7404 53524 7410
rect 53472 7346 53524 7352
rect 53380 7200 53432 7206
rect 53380 7142 53432 7148
rect 53392 7041 53420 7142
rect 53378 7032 53434 7041
rect 53378 6967 53434 6976
rect 53288 6724 53340 6730
rect 53288 6666 53340 6672
rect 53300 6458 53328 6666
rect 53288 6452 53340 6458
rect 53288 6394 53340 6400
rect 53104 6316 53156 6322
rect 53104 6258 53156 6264
rect 52920 6248 52972 6254
rect 52920 6190 52972 6196
rect 53012 6248 53064 6254
rect 53012 6190 53064 6196
rect 52932 5914 52960 6190
rect 52920 5908 52972 5914
rect 52920 5850 52972 5856
rect 52932 5574 52960 5850
rect 53116 5778 53144 6258
rect 53472 6112 53524 6118
rect 53472 6054 53524 6060
rect 53104 5772 53156 5778
rect 53104 5714 53156 5720
rect 53484 5710 53512 6054
rect 53576 5914 53604 10950
rect 53668 10033 53696 12135
rect 53760 11218 53788 12718
rect 53840 12232 53892 12238
rect 53840 12174 53892 12180
rect 53748 11212 53800 11218
rect 53748 11154 53800 11160
rect 53748 10260 53800 10266
rect 53748 10202 53800 10208
rect 53760 10062 53788 10202
rect 53748 10056 53800 10062
rect 53654 10024 53710 10033
rect 53748 9998 53800 10004
rect 53852 9994 53880 12174
rect 53654 9959 53710 9968
rect 53840 9988 53892 9994
rect 53668 9586 53696 9959
rect 53840 9930 53892 9936
rect 53748 9920 53800 9926
rect 53748 9862 53800 9868
rect 53760 9625 53788 9862
rect 53746 9616 53802 9625
rect 53656 9580 53708 9586
rect 53746 9551 53802 9560
rect 53656 9522 53708 9528
rect 53748 9512 53800 9518
rect 53748 9454 53800 9460
rect 53656 7812 53708 7818
rect 53656 7754 53708 7760
rect 53668 7206 53696 7754
rect 53656 7200 53708 7206
rect 53656 7142 53708 7148
rect 53564 5908 53616 5914
rect 53564 5850 53616 5856
rect 53472 5704 53524 5710
rect 53472 5646 53524 5652
rect 52920 5568 52972 5574
rect 52920 5510 52972 5516
rect 53484 5234 53512 5646
rect 53760 5302 53788 9454
rect 53944 9042 53972 13806
rect 54036 12442 54064 14962
rect 54116 14884 54168 14890
rect 54116 14826 54168 14832
rect 54024 12436 54076 12442
rect 54024 12378 54076 12384
rect 54128 11762 54156 14826
rect 54208 13932 54260 13938
rect 54208 13874 54260 13880
rect 54220 13462 54248 13874
rect 54208 13456 54260 13462
rect 54208 13398 54260 13404
rect 54208 13252 54260 13258
rect 54208 13194 54260 13200
rect 54220 12481 54248 13194
rect 54206 12472 54262 12481
rect 54206 12407 54262 12416
rect 54208 12096 54260 12102
rect 54208 12038 54260 12044
rect 54220 11898 54248 12038
rect 54208 11892 54260 11898
rect 54208 11834 54260 11840
rect 54116 11756 54168 11762
rect 54116 11698 54168 11704
rect 54208 11688 54260 11694
rect 54208 11630 54260 11636
rect 54220 11354 54248 11630
rect 54312 11354 54340 16487
rect 54484 16458 54536 16464
rect 54496 16250 54524 16458
rect 54484 16244 54536 16250
rect 54484 16186 54536 16192
rect 54496 15978 54524 16186
rect 54484 15972 54536 15978
rect 54484 15914 54536 15920
rect 54484 15428 54536 15434
rect 54484 15370 54536 15376
rect 54392 15020 54444 15026
rect 54392 14962 54444 14968
rect 54404 14618 54432 14962
rect 54392 14612 54444 14618
rect 54392 14554 54444 14560
rect 54392 14272 54444 14278
rect 54392 14214 54444 14220
rect 54404 13530 54432 14214
rect 54392 13524 54444 13530
rect 54392 13466 54444 13472
rect 54392 12708 54444 12714
rect 54496 12696 54524 15370
rect 54588 15162 54616 17190
rect 54668 16584 54720 16590
rect 54668 16526 54720 16532
rect 54576 15156 54628 15162
rect 54576 15098 54628 15104
rect 54680 15094 54708 16526
rect 54772 15960 54800 18022
rect 55600 17882 55628 22578
rect 55692 22438 55720 23054
rect 55864 22568 55916 22574
rect 55864 22510 55916 22516
rect 55680 22432 55732 22438
rect 55680 22374 55732 22380
rect 55876 22098 55904 22510
rect 55864 22092 55916 22098
rect 55864 22034 55916 22040
rect 55680 20936 55732 20942
rect 55680 20878 55732 20884
rect 55692 20262 55720 20878
rect 55680 20256 55732 20262
rect 55680 20198 55732 20204
rect 56336 20058 56364 23582
rect 56876 23530 56928 23536
rect 56968 23044 57020 23050
rect 56968 22986 57020 22992
rect 56980 22778 57008 22986
rect 56968 22772 57020 22778
rect 56968 22714 57020 22720
rect 56600 22704 56652 22710
rect 56600 22646 56652 22652
rect 56784 22704 56836 22710
rect 56784 22646 56836 22652
rect 56508 22432 56560 22438
rect 56508 22374 56560 22380
rect 56520 22030 56548 22374
rect 56508 22024 56560 22030
rect 56508 21966 56560 21972
rect 56612 21894 56640 22646
rect 56796 21962 56824 22646
rect 56784 21956 56836 21962
rect 56784 21898 56836 21904
rect 56600 21888 56652 21894
rect 56600 21830 56652 21836
rect 56796 21690 56824 21898
rect 56784 21684 56836 21690
rect 56784 21626 56836 21632
rect 56876 21548 56928 21554
rect 56876 21490 56928 21496
rect 56968 21548 57020 21554
rect 56968 21490 57020 21496
rect 56888 21146 56916 21490
rect 56980 21146 57008 21490
rect 56876 21140 56928 21146
rect 56876 21082 56928 21088
rect 56968 21140 57020 21146
rect 56968 21082 57020 21088
rect 56508 20868 56560 20874
rect 56508 20810 56560 20816
rect 56520 20398 56548 20810
rect 56600 20800 56652 20806
rect 56600 20742 56652 20748
rect 56612 20466 56640 20742
rect 56980 20534 57008 21082
rect 56968 20528 57020 20534
rect 56968 20470 57020 20476
rect 56600 20460 56652 20466
rect 56600 20402 56652 20408
rect 56508 20392 56560 20398
rect 56508 20334 56560 20340
rect 56324 20052 56376 20058
rect 56324 19994 56376 20000
rect 56520 19854 56548 20334
rect 56692 20256 56744 20262
rect 56692 20198 56744 20204
rect 56600 19916 56652 19922
rect 56600 19858 56652 19864
rect 56508 19848 56560 19854
rect 56428 19796 56508 19802
rect 56428 19790 56560 19796
rect 56428 19774 56548 19790
rect 56428 19718 56456 19774
rect 56416 19712 56468 19718
rect 56416 19654 56468 19660
rect 56048 19440 56100 19446
rect 56048 19382 56100 19388
rect 55956 19304 56008 19310
rect 55956 19246 56008 19252
rect 55772 18828 55824 18834
rect 55772 18770 55824 18776
rect 55680 18624 55732 18630
rect 55680 18566 55732 18572
rect 55692 18358 55720 18566
rect 55680 18352 55732 18358
rect 55680 18294 55732 18300
rect 55588 17876 55640 17882
rect 55588 17818 55640 17824
rect 55692 17746 55720 18294
rect 55784 18290 55812 18770
rect 55968 18698 55996 19246
rect 55956 18692 56008 18698
rect 55956 18634 56008 18640
rect 55968 18290 55996 18634
rect 56060 18630 56088 19382
rect 56428 19378 56456 19654
rect 56416 19372 56468 19378
rect 56416 19314 56468 19320
rect 56048 18624 56100 18630
rect 56048 18566 56100 18572
rect 55772 18284 55824 18290
rect 55772 18226 55824 18232
rect 55956 18284 56008 18290
rect 55956 18226 56008 18232
rect 55968 17864 55996 18226
rect 55876 17836 55996 17864
rect 55680 17740 55732 17746
rect 55680 17682 55732 17688
rect 55876 17678 55904 17836
rect 55956 17740 56008 17746
rect 55956 17682 56008 17688
rect 55864 17672 55916 17678
rect 55864 17614 55916 17620
rect 54944 17536 54996 17542
rect 54944 17478 54996 17484
rect 54852 17196 54904 17202
rect 54852 17138 54904 17144
rect 54864 16794 54892 17138
rect 54852 16788 54904 16794
rect 54852 16730 54904 16736
rect 54852 15972 54904 15978
rect 54772 15932 54852 15960
rect 54852 15914 54904 15920
rect 54668 15088 54720 15094
rect 54668 15030 54720 15036
rect 54576 14408 54628 14414
rect 54576 14350 54628 14356
rect 54588 13938 54616 14350
rect 54680 14074 54708 15030
rect 54864 14278 54892 15914
rect 54956 15706 54984 17478
rect 55876 17202 55904 17614
rect 55968 17202 55996 17682
rect 55864 17196 55916 17202
rect 55864 17138 55916 17144
rect 55956 17196 56008 17202
rect 55956 17138 56008 17144
rect 55680 17060 55732 17066
rect 55680 17002 55732 17008
rect 55496 16992 55548 16998
rect 55496 16934 55548 16940
rect 55508 16590 55536 16934
rect 55036 16584 55088 16590
rect 55036 16526 55088 16532
rect 55496 16584 55548 16590
rect 55496 16526 55548 16532
rect 55588 16584 55640 16590
rect 55588 16526 55640 16532
rect 54944 15700 54996 15706
rect 54944 15642 54996 15648
rect 54852 14272 54904 14278
rect 54852 14214 54904 14220
rect 54668 14068 54720 14074
rect 54668 14010 54720 14016
rect 54852 14000 54904 14006
rect 54852 13942 54904 13948
rect 54576 13932 54628 13938
rect 54576 13874 54628 13880
rect 54588 13530 54616 13874
rect 54576 13524 54628 13530
rect 54576 13466 54628 13472
rect 54864 12850 54892 13942
rect 55048 12850 55076 16526
rect 55220 16108 55272 16114
rect 55220 16050 55272 16056
rect 55128 15904 55180 15910
rect 55128 15846 55180 15852
rect 55140 14618 55168 15846
rect 55232 15502 55260 16050
rect 55508 16046 55536 16526
rect 55600 16114 55628 16526
rect 55692 16250 55720 17002
rect 56060 16794 56088 18566
rect 56428 17338 56456 19314
rect 56612 19310 56640 19858
rect 56600 19304 56652 19310
rect 56600 19246 56652 19252
rect 56600 17740 56652 17746
rect 56600 17682 56652 17688
rect 56416 17332 56468 17338
rect 56416 17274 56468 17280
rect 56508 17196 56560 17202
rect 56508 17138 56560 17144
rect 56048 16788 56100 16794
rect 56048 16730 56100 16736
rect 56520 16658 56548 17138
rect 56612 16794 56640 17682
rect 56600 16788 56652 16794
rect 56600 16730 56652 16736
rect 56508 16652 56560 16658
rect 56508 16594 56560 16600
rect 56520 16250 56548 16594
rect 56704 16522 56732 20198
rect 56784 16584 56836 16590
rect 56784 16526 56836 16532
rect 56692 16516 56744 16522
rect 56692 16458 56744 16464
rect 56600 16448 56652 16454
rect 56600 16390 56652 16396
rect 55680 16244 55732 16250
rect 55680 16186 55732 16192
rect 56508 16244 56560 16250
rect 56508 16186 56560 16192
rect 55588 16108 55640 16114
rect 55588 16050 55640 16056
rect 55496 16040 55548 16046
rect 55496 15982 55548 15988
rect 55220 15496 55272 15502
rect 55220 15438 55272 15444
rect 55218 15192 55274 15201
rect 55218 15127 55274 15136
rect 55232 15026 55260 15127
rect 55508 15026 55536 15982
rect 55600 15745 55628 16050
rect 55586 15736 55642 15745
rect 55586 15671 55642 15680
rect 55600 15026 55628 15671
rect 55220 15020 55272 15026
rect 55496 15020 55548 15026
rect 55272 14980 55444 15008
rect 55220 14962 55272 14968
rect 55128 14612 55180 14618
rect 55128 14554 55180 14560
rect 55140 14074 55168 14554
rect 55218 14512 55274 14521
rect 55218 14447 55274 14456
rect 55232 14074 55260 14447
rect 55128 14068 55180 14074
rect 55128 14010 55180 14016
rect 55220 14068 55272 14074
rect 55220 14010 55272 14016
rect 55128 13456 55180 13462
rect 55128 13398 55180 13404
rect 54852 12844 54904 12850
rect 54852 12786 54904 12792
rect 55036 12844 55088 12850
rect 55036 12786 55088 12792
rect 54444 12668 54524 12696
rect 54392 12650 54444 12656
rect 54208 11348 54260 11354
rect 54208 11290 54260 11296
rect 54300 11348 54352 11354
rect 54300 11290 54352 11296
rect 54404 11200 54432 12650
rect 54758 12472 54814 12481
rect 54758 12407 54814 12416
rect 54484 12368 54536 12374
rect 54484 12310 54536 12316
rect 54496 11830 54524 12310
rect 54668 12232 54720 12238
rect 54668 12174 54720 12180
rect 54484 11824 54536 11830
rect 54484 11766 54536 11772
rect 54576 11756 54628 11762
rect 54576 11698 54628 11704
rect 54220 11172 54432 11200
rect 54484 11212 54536 11218
rect 54116 11144 54168 11150
rect 54116 11086 54168 11092
rect 54022 10840 54078 10849
rect 54022 10775 54024 10784
rect 54076 10775 54078 10784
rect 54024 10746 54076 10752
rect 54128 10266 54156 11086
rect 54220 10810 54248 11172
rect 54484 11154 54536 11160
rect 54392 11076 54444 11082
rect 54392 11018 54444 11024
rect 54298 10976 54354 10985
rect 54298 10911 54354 10920
rect 54208 10804 54260 10810
rect 54208 10746 54260 10752
rect 54312 10674 54340 10911
rect 54208 10668 54260 10674
rect 54208 10610 54260 10616
rect 54300 10668 54352 10674
rect 54300 10610 54352 10616
rect 54116 10260 54168 10266
rect 54116 10202 54168 10208
rect 54024 9376 54076 9382
rect 54024 9318 54076 9324
rect 54036 9042 54064 9318
rect 54220 9178 54248 10610
rect 54208 9172 54260 9178
rect 54208 9114 54260 9120
rect 53932 9036 53984 9042
rect 53932 8978 53984 8984
rect 54024 9036 54076 9042
rect 54024 8978 54076 8984
rect 53944 7970 53972 8978
rect 54404 8974 54432 11018
rect 54496 10606 54524 11154
rect 54588 10674 54616 11698
rect 54576 10668 54628 10674
rect 54576 10610 54628 10616
rect 54484 10600 54536 10606
rect 54484 10542 54536 10548
rect 54680 10441 54708 12174
rect 54666 10432 54722 10441
rect 54666 10367 54722 10376
rect 54576 9512 54628 9518
rect 54576 9454 54628 9460
rect 54484 9104 54536 9110
rect 54484 9046 54536 9052
rect 54392 8968 54444 8974
rect 54392 8910 54444 8916
rect 54024 8628 54076 8634
rect 54024 8570 54076 8576
rect 54036 8430 54064 8570
rect 54024 8424 54076 8430
rect 54024 8366 54076 8372
rect 53852 7942 53972 7970
rect 53852 6186 53880 7942
rect 53932 7540 53984 7546
rect 53932 7482 53984 7488
rect 53944 7410 53972 7482
rect 53932 7404 53984 7410
rect 53932 7346 53984 7352
rect 53840 6180 53892 6186
rect 53840 6122 53892 6128
rect 53748 5296 53800 5302
rect 53748 5238 53800 5244
rect 53472 5228 53524 5234
rect 53472 5170 53524 5176
rect 52828 4820 52880 4826
rect 52828 4762 52880 4768
rect 53104 4752 53156 4758
rect 53104 4694 53156 4700
rect 53116 4214 53144 4694
rect 52552 4208 52604 4214
rect 52552 4150 52604 4156
rect 53104 4208 53156 4214
rect 53104 4150 53156 4156
rect 53484 3942 53512 5170
rect 54036 4826 54064 8366
rect 54300 8356 54352 8362
rect 54300 8298 54352 8304
rect 54206 8256 54262 8265
rect 54206 8191 54262 8200
rect 54116 7880 54168 7886
rect 54116 7822 54168 7828
rect 54128 7478 54156 7822
rect 54220 7546 54248 8191
rect 54208 7540 54260 7546
rect 54208 7482 54260 7488
rect 54116 7472 54168 7478
rect 54116 7414 54168 7420
rect 54312 7342 54340 8298
rect 54404 8294 54432 8910
rect 54392 8288 54444 8294
rect 54392 8230 54444 8236
rect 54404 7886 54432 8230
rect 54392 7880 54444 7886
rect 54392 7822 54444 7828
rect 54496 7410 54524 9046
rect 54588 8838 54616 9454
rect 54576 8832 54628 8838
rect 54576 8774 54628 8780
rect 54588 8566 54616 8774
rect 54680 8634 54708 10367
rect 54668 8628 54720 8634
rect 54668 8570 54720 8576
rect 54576 8560 54628 8566
rect 54576 8502 54628 8508
rect 54772 8022 54800 12407
rect 54864 12102 54892 12786
rect 54944 12776 54996 12782
rect 54944 12718 54996 12724
rect 54956 12442 54984 12718
rect 54944 12436 54996 12442
rect 54944 12378 54996 12384
rect 54852 12096 54904 12102
rect 54852 12038 54904 12044
rect 54852 11620 54904 11626
rect 54852 11562 54904 11568
rect 54864 11200 54892 11562
rect 54956 11268 54984 12378
rect 55048 11762 55076 12786
rect 55036 11756 55088 11762
rect 55036 11698 55088 11704
rect 54956 11240 55076 11268
rect 54864 11172 54984 11200
rect 54852 11076 54904 11082
rect 54852 11018 54904 11024
rect 54864 9382 54892 11018
rect 54852 9376 54904 9382
rect 54852 9318 54904 9324
rect 54864 8634 54892 9318
rect 54852 8628 54904 8634
rect 54852 8570 54904 8576
rect 54852 8492 54904 8498
rect 54852 8434 54904 8440
rect 54760 8016 54812 8022
rect 54760 7958 54812 7964
rect 54864 7954 54892 8434
rect 54852 7948 54904 7954
rect 54852 7890 54904 7896
rect 54760 7880 54812 7886
rect 54760 7822 54812 7828
rect 54484 7404 54536 7410
rect 54484 7346 54536 7352
rect 54668 7404 54720 7410
rect 54668 7346 54720 7352
rect 54300 7336 54352 7342
rect 54300 7278 54352 7284
rect 54680 6934 54708 7346
rect 54772 7206 54800 7822
rect 54864 7410 54892 7890
rect 54852 7404 54904 7410
rect 54852 7346 54904 7352
rect 54760 7200 54812 7206
rect 54760 7142 54812 7148
rect 54668 6928 54720 6934
rect 54668 6870 54720 6876
rect 54772 6798 54800 7142
rect 54760 6792 54812 6798
rect 54760 6734 54812 6740
rect 54850 6760 54906 6769
rect 54116 6656 54168 6662
rect 54116 6598 54168 6604
rect 54208 6656 54260 6662
rect 54208 6598 54260 6604
rect 54128 6118 54156 6598
rect 54220 6254 54248 6598
rect 54208 6248 54260 6254
rect 54208 6190 54260 6196
rect 54116 6112 54168 6118
rect 54116 6054 54168 6060
rect 54116 5772 54168 5778
rect 54116 5714 54168 5720
rect 54128 5370 54156 5714
rect 54220 5710 54248 6190
rect 54772 5778 54800 6734
rect 54850 6695 54852 6704
rect 54904 6695 54906 6704
rect 54852 6666 54904 6672
rect 54852 6452 54904 6458
rect 54852 6394 54904 6400
rect 54760 5772 54812 5778
rect 54760 5714 54812 5720
rect 54864 5710 54892 6394
rect 54208 5704 54260 5710
rect 54208 5646 54260 5652
rect 54852 5704 54904 5710
rect 54852 5646 54904 5652
rect 54116 5364 54168 5370
rect 54116 5306 54168 5312
rect 54024 4820 54076 4826
rect 54024 4762 54076 4768
rect 54220 4690 54248 5646
rect 54852 5568 54904 5574
rect 54852 5510 54904 5516
rect 54864 5370 54892 5510
rect 54852 5364 54904 5370
rect 54852 5306 54904 5312
rect 54668 5160 54720 5166
rect 54668 5102 54720 5108
rect 54208 4684 54260 4690
rect 54208 4626 54260 4632
rect 54220 4282 54248 4626
rect 54576 4616 54628 4622
rect 54576 4558 54628 4564
rect 54208 4276 54260 4282
rect 54208 4218 54260 4224
rect 54220 4078 54248 4218
rect 54208 4072 54260 4078
rect 54208 4014 54260 4020
rect 53472 3936 53524 3942
rect 53472 3878 53524 3884
rect 52276 3528 52328 3534
rect 52276 3470 52328 3476
rect 52288 3194 52316 3470
rect 53484 3398 53512 3878
rect 54220 3738 54248 4014
rect 54208 3732 54260 3738
rect 54208 3674 54260 3680
rect 53472 3392 53524 3398
rect 53472 3334 53524 3340
rect 53484 3194 53512 3334
rect 54220 3194 54248 3674
rect 54588 3194 54616 4558
rect 54680 4010 54708 5102
rect 54956 4214 54984 11172
rect 55048 11150 55076 11240
rect 55036 11144 55088 11150
rect 55036 11086 55088 11092
rect 55140 10849 55168 13398
rect 55416 13308 55444 14980
rect 55496 14962 55548 14968
rect 55588 15020 55640 15026
rect 55588 14962 55640 14968
rect 55508 14006 55536 14962
rect 55496 14000 55548 14006
rect 55496 13942 55548 13948
rect 55600 13462 55628 14962
rect 55692 14890 55720 16186
rect 56612 15910 56640 16390
rect 56600 15904 56652 15910
rect 56600 15846 56652 15852
rect 56612 15570 56640 15846
rect 56796 15638 56824 16526
rect 56968 16516 57020 16522
rect 56968 16458 57020 16464
rect 56784 15632 56836 15638
rect 56784 15574 56836 15580
rect 56600 15564 56652 15570
rect 56600 15506 56652 15512
rect 56692 15496 56744 15502
rect 56692 15438 56744 15444
rect 56232 15360 56284 15366
rect 56232 15302 56284 15308
rect 55956 15020 56008 15026
rect 55956 14962 56008 14968
rect 55680 14884 55732 14890
rect 55680 14826 55732 14832
rect 55692 14414 55720 14826
rect 55680 14408 55732 14414
rect 55680 14350 55732 14356
rect 55588 13456 55640 13462
rect 55588 13398 55640 13404
rect 55416 13280 55628 13308
rect 55404 12640 55456 12646
rect 55402 12608 55404 12617
rect 55456 12608 55458 12617
rect 55402 12543 55458 12552
rect 55220 12232 55272 12238
rect 55220 12174 55272 12180
rect 55126 10840 55182 10849
rect 55126 10775 55128 10784
rect 55180 10775 55182 10784
rect 55128 10746 55180 10752
rect 55140 10715 55168 10746
rect 55128 8016 55180 8022
rect 55128 7958 55180 7964
rect 55036 6724 55088 6730
rect 55036 6666 55088 6672
rect 55048 5778 55076 6666
rect 55140 6390 55168 7958
rect 55232 7449 55260 12174
rect 55312 12096 55364 12102
rect 55312 12038 55364 12044
rect 55324 11082 55352 12038
rect 55312 11076 55364 11082
rect 55312 11018 55364 11024
rect 55312 10464 55364 10470
rect 55312 10406 55364 10412
rect 55324 9926 55352 10406
rect 55312 9920 55364 9926
rect 55312 9862 55364 9868
rect 55416 9042 55444 12543
rect 55496 12368 55548 12374
rect 55494 12336 55496 12345
rect 55548 12336 55550 12345
rect 55494 12271 55550 12280
rect 55496 12164 55548 12170
rect 55496 12106 55548 12112
rect 55508 11830 55536 12106
rect 55496 11824 55548 11830
rect 55496 11766 55548 11772
rect 55508 10742 55536 11766
rect 55496 10736 55548 10742
rect 55496 10678 55548 10684
rect 55496 9444 55548 9450
rect 55496 9386 55548 9392
rect 55404 9036 55456 9042
rect 55404 8978 55456 8984
rect 55312 8628 55364 8634
rect 55312 8570 55364 8576
rect 55218 7440 55274 7449
rect 55218 7375 55274 7384
rect 55232 6866 55260 7375
rect 55220 6860 55272 6866
rect 55220 6802 55272 6808
rect 55128 6384 55180 6390
rect 55128 6326 55180 6332
rect 55036 5772 55088 5778
rect 55036 5714 55088 5720
rect 55048 5030 55076 5714
rect 55140 5642 55168 6326
rect 55128 5636 55180 5642
rect 55128 5578 55180 5584
rect 55140 5302 55168 5578
rect 55324 5370 55352 8570
rect 55416 8362 55444 8978
rect 55508 8498 55536 9386
rect 55496 8492 55548 8498
rect 55496 8434 55548 8440
rect 55404 8356 55456 8362
rect 55404 8298 55456 8304
rect 55496 7200 55548 7206
rect 55496 7142 55548 7148
rect 55508 5846 55536 7142
rect 55496 5840 55548 5846
rect 55496 5782 55548 5788
rect 55312 5364 55364 5370
rect 55312 5306 55364 5312
rect 55128 5296 55180 5302
rect 55128 5238 55180 5244
rect 55036 5024 55088 5030
rect 55036 4966 55088 4972
rect 55140 4282 55168 5238
rect 55220 4752 55272 4758
rect 55220 4694 55272 4700
rect 55128 4276 55180 4282
rect 55128 4218 55180 4224
rect 54944 4208 54996 4214
rect 54944 4150 54996 4156
rect 54668 4004 54720 4010
rect 54668 3946 54720 3952
rect 54680 3738 54708 3946
rect 54668 3732 54720 3738
rect 54668 3674 54720 3680
rect 55232 3194 55260 4694
rect 55600 4622 55628 13280
rect 55864 13184 55916 13190
rect 55968 13138 55996 14962
rect 56244 14618 56272 15302
rect 56232 14612 56284 14618
rect 56232 14554 56284 14560
rect 56704 14278 56732 15438
rect 56980 15026 57008 16458
rect 56968 15020 57020 15026
rect 56968 14962 57020 14968
rect 56692 14272 56744 14278
rect 56692 14214 56744 14220
rect 56232 14068 56284 14074
rect 56232 14010 56284 14016
rect 56048 13932 56100 13938
rect 56048 13874 56100 13880
rect 56060 13258 56088 13874
rect 56244 13326 56272 14010
rect 56416 13932 56468 13938
rect 56416 13874 56468 13880
rect 56428 13462 56456 13874
rect 56508 13864 56560 13870
rect 56508 13806 56560 13812
rect 56520 13530 56548 13806
rect 56598 13560 56654 13569
rect 56508 13524 56560 13530
rect 56598 13495 56600 13504
rect 56508 13466 56560 13472
rect 56652 13495 56654 13504
rect 56600 13466 56652 13472
rect 56416 13456 56468 13462
rect 56416 13398 56468 13404
rect 56232 13320 56284 13326
rect 56232 13262 56284 13268
rect 56048 13252 56100 13258
rect 56048 13194 56100 13200
rect 55916 13132 55996 13138
rect 55864 13126 55996 13132
rect 55876 13110 55996 13126
rect 55772 12776 55824 12782
rect 55772 12718 55824 12724
rect 55680 12640 55732 12646
rect 55680 12582 55732 12588
rect 55692 12238 55720 12582
rect 55680 12232 55732 12238
rect 55680 12174 55732 12180
rect 55680 12096 55732 12102
rect 55784 12084 55812 12718
rect 55732 12056 55812 12084
rect 55680 12038 55732 12044
rect 55692 11898 55720 12038
rect 55680 11892 55732 11898
rect 55680 11834 55732 11840
rect 55772 11824 55824 11830
rect 55772 11766 55824 11772
rect 55680 11552 55732 11558
rect 55680 11494 55732 11500
rect 55692 11200 55720 11494
rect 55784 11354 55812 11766
rect 55772 11348 55824 11354
rect 55772 11290 55824 11296
rect 55692 11172 55812 11200
rect 55680 11076 55732 11082
rect 55680 11018 55732 11024
rect 55692 10198 55720 11018
rect 55784 11014 55812 11172
rect 55772 11008 55824 11014
rect 55772 10950 55824 10956
rect 55680 10192 55732 10198
rect 55680 10134 55732 10140
rect 55692 9178 55720 10134
rect 55680 9172 55732 9178
rect 55680 9114 55732 9120
rect 55692 7750 55720 9114
rect 55876 8106 55904 13110
rect 55956 12300 56008 12306
rect 55956 12242 56008 12248
rect 55968 11898 55996 12242
rect 55956 11892 56008 11898
rect 55956 11834 56008 11840
rect 56060 9654 56088 13194
rect 56232 13184 56284 13190
rect 56232 13126 56284 13132
rect 56244 12918 56272 13126
rect 56232 12912 56284 12918
rect 56232 12854 56284 12860
rect 56324 10736 56376 10742
rect 56244 10696 56324 10724
rect 56140 10668 56192 10674
rect 56140 10610 56192 10616
rect 56152 10062 56180 10610
rect 56140 10056 56192 10062
rect 56140 9998 56192 10004
rect 56152 9722 56180 9998
rect 56140 9716 56192 9722
rect 56140 9658 56192 9664
rect 56048 9648 56100 9654
rect 56048 9590 56100 9596
rect 56060 8498 56088 9590
rect 56048 8492 56100 8498
rect 56100 8452 56180 8480
rect 56048 8434 56100 8440
rect 55876 8090 56088 8106
rect 55876 8084 56100 8090
rect 55876 8078 56048 8084
rect 56048 8026 56100 8032
rect 55864 8016 55916 8022
rect 55864 7958 55916 7964
rect 55876 7886 55904 7958
rect 56152 7954 56180 8452
rect 56140 7948 56192 7954
rect 56140 7890 56192 7896
rect 55864 7880 55916 7886
rect 55864 7822 55916 7828
rect 55680 7744 55732 7750
rect 55680 7686 55732 7692
rect 55692 7206 55720 7686
rect 56152 7478 56180 7890
rect 56140 7472 56192 7478
rect 56140 7414 56192 7420
rect 55680 7200 55732 7206
rect 55680 7142 55732 7148
rect 56244 6866 56272 10696
rect 56324 10678 56376 10684
rect 56428 10062 56456 13398
rect 56520 11014 56548 13466
rect 56704 12646 56732 14214
rect 56968 12912 57020 12918
rect 56968 12854 57020 12860
rect 56980 12714 57008 12854
rect 56968 12708 57020 12714
rect 56968 12650 57020 12656
rect 56692 12640 56744 12646
rect 56692 12582 56744 12588
rect 56508 11008 56560 11014
rect 56508 10950 56560 10956
rect 56692 11008 56744 11014
rect 56692 10950 56744 10956
rect 56416 10056 56468 10062
rect 56416 9998 56468 10004
rect 56428 9738 56456 9998
rect 56336 9722 56456 9738
rect 56336 9716 56468 9722
rect 56336 9710 56416 9716
rect 56336 9110 56364 9710
rect 56416 9658 56468 9664
rect 56416 9580 56468 9586
rect 56416 9522 56468 9528
rect 56324 9104 56376 9110
rect 56324 9046 56376 9052
rect 56428 8945 56456 9522
rect 56520 8974 56548 10950
rect 56598 10704 56654 10713
rect 56598 10639 56654 10648
rect 56612 9178 56640 10639
rect 56704 10266 56732 10950
rect 56784 10464 56836 10470
rect 56784 10406 56836 10412
rect 56692 10260 56744 10266
rect 56692 10202 56744 10208
rect 56600 9172 56652 9178
rect 56600 9114 56652 9120
rect 56508 8968 56560 8974
rect 56414 8936 56470 8945
rect 56508 8910 56560 8916
rect 56414 8871 56470 8880
rect 56428 8498 56456 8871
rect 56416 8492 56468 8498
rect 56416 8434 56468 8440
rect 56324 7200 56376 7206
rect 56324 7142 56376 7148
rect 56336 7002 56364 7142
rect 56324 6996 56376 7002
rect 56324 6938 56376 6944
rect 56232 6860 56284 6866
rect 56232 6802 56284 6808
rect 56520 6186 56548 8910
rect 56704 8838 56732 10202
rect 56796 10130 56824 10406
rect 56784 10124 56836 10130
rect 56784 10066 56836 10072
rect 56980 9926 57008 12650
rect 56968 9920 57020 9926
rect 56968 9862 57020 9868
rect 56876 9648 56928 9654
rect 56876 9590 56928 9596
rect 56888 9450 56916 9590
rect 56876 9444 56928 9450
rect 56876 9386 56928 9392
rect 56784 9376 56836 9382
rect 56784 9318 56836 9324
rect 56692 8832 56744 8838
rect 56692 8774 56744 8780
rect 56704 8634 56732 8774
rect 56692 8628 56744 8634
rect 56692 8570 56744 8576
rect 56796 7886 56824 9318
rect 56888 8838 56916 9386
rect 56876 8832 56928 8838
rect 56876 8774 56928 8780
rect 56784 7880 56836 7886
rect 56784 7822 56836 7828
rect 56796 7546 56824 7822
rect 56784 7540 56836 7546
rect 56784 7482 56836 7488
rect 56508 6180 56560 6186
rect 56508 6122 56560 6128
rect 56520 5914 56548 6122
rect 56888 6118 56916 8774
rect 56980 7274 57008 9862
rect 56968 7268 57020 7274
rect 56968 7210 57020 7216
rect 56600 6112 56652 6118
rect 56600 6054 56652 6060
rect 56876 6112 56928 6118
rect 56876 6054 56928 6060
rect 56508 5908 56560 5914
rect 56508 5850 56560 5856
rect 56048 5228 56100 5234
rect 56048 5170 56100 5176
rect 56060 4826 56088 5170
rect 56508 5024 56560 5030
rect 56612 5012 56640 6054
rect 56560 4984 56640 5012
rect 56508 4966 56560 4972
rect 56048 4820 56100 4826
rect 56048 4762 56100 4768
rect 55588 4616 55640 4622
rect 55588 4558 55640 4564
rect 55496 4208 55548 4214
rect 55496 4150 55548 4156
rect 55508 3738 55536 4150
rect 55496 3732 55548 3738
rect 55496 3674 55548 3680
rect 56520 3670 56548 4966
rect 56508 3664 56560 3670
rect 56508 3606 56560 3612
rect 52276 3188 52328 3194
rect 52276 3130 52328 3136
rect 53472 3188 53524 3194
rect 53472 3130 53524 3136
rect 54208 3188 54260 3194
rect 54208 3130 54260 3136
rect 54576 3188 54628 3194
rect 54576 3130 54628 3136
rect 55220 3188 55272 3194
rect 55220 3130 55272 3136
rect 52184 3052 52236 3058
rect 52184 2994 52236 3000
rect 53484 2650 53512 3130
rect 57072 2774 57100 25162
rect 57244 18624 57296 18630
rect 57244 18566 57296 18572
rect 57256 17542 57284 18566
rect 57244 17536 57296 17542
rect 57244 17478 57296 17484
rect 57152 15904 57204 15910
rect 57152 15846 57204 15852
rect 57164 15434 57192 15846
rect 57152 15428 57204 15434
rect 57152 15370 57204 15376
rect 57348 14006 57376 54470
rect 57520 42560 57572 42566
rect 57520 42502 57572 42508
rect 57532 29782 57560 42502
rect 57520 29776 57572 29782
rect 57520 29718 57572 29724
rect 57520 26784 57572 26790
rect 57520 26726 57572 26732
rect 57428 26512 57480 26518
rect 57428 26454 57480 26460
rect 57440 25906 57468 26454
rect 57428 25900 57480 25906
rect 57428 25842 57480 25848
rect 57532 25294 57560 26726
rect 57612 25900 57664 25906
rect 57612 25842 57664 25848
rect 57624 25430 57652 25842
rect 57612 25424 57664 25430
rect 57612 25366 57664 25372
rect 57520 25288 57572 25294
rect 57520 25230 57572 25236
rect 57428 23656 57480 23662
rect 57428 23598 57480 23604
rect 57440 23050 57468 23598
rect 57624 23322 57652 25366
rect 57612 23316 57664 23322
rect 57612 23258 57664 23264
rect 57428 23044 57480 23050
rect 57428 22986 57480 22992
rect 57440 22234 57468 22986
rect 57428 22228 57480 22234
rect 57428 22170 57480 22176
rect 57716 22094 57744 57190
rect 58256 54528 58308 54534
rect 58254 54496 58256 54505
rect 58308 54496 58310 54505
rect 58254 54431 58310 54440
rect 57796 48748 57848 48754
rect 57796 48690 57848 48696
rect 57808 48550 57836 48690
rect 57796 48544 57848 48550
rect 57796 48486 57848 48492
rect 58256 48544 58308 48550
rect 58256 48486 58308 48492
rect 57808 25498 57836 48486
rect 58268 48385 58296 48486
rect 58254 48376 58310 48385
rect 58254 48311 58310 48320
rect 58256 42560 58308 42566
rect 58256 42502 58308 42508
rect 58268 42265 58296 42502
rect 58254 42256 58310 42265
rect 58254 42191 58310 42200
rect 57980 37256 58032 37262
rect 57980 37198 58032 37204
rect 57992 35894 58020 37198
rect 58256 37120 58308 37126
rect 58256 37062 58308 37068
rect 58268 36825 58296 37062
rect 58254 36816 58310 36825
rect 58254 36751 58310 36760
rect 57992 35866 58112 35894
rect 57888 27464 57940 27470
rect 57888 27406 57940 27412
rect 57900 26450 57928 27406
rect 57888 26444 57940 26450
rect 57888 26386 57940 26392
rect 57796 25492 57848 25498
rect 57796 25434 57848 25440
rect 58084 24410 58112 35866
rect 58164 30728 58216 30734
rect 58164 30670 58216 30676
rect 58254 30696 58310 30705
rect 58072 24404 58124 24410
rect 58072 24346 58124 24352
rect 57888 24200 57940 24206
rect 57888 24142 57940 24148
rect 58072 24200 58124 24206
rect 58072 24142 58124 24148
rect 57796 23520 57848 23526
rect 57796 23462 57848 23468
rect 57808 22098 57836 23462
rect 57624 22066 57744 22094
rect 57796 22092 57848 22098
rect 57520 20868 57572 20874
rect 57520 20810 57572 20816
rect 57532 20602 57560 20810
rect 57520 20596 57572 20602
rect 57520 20538 57572 20544
rect 57428 19916 57480 19922
rect 57428 19858 57480 19864
rect 57440 19514 57468 19858
rect 57428 19508 57480 19514
rect 57428 19450 57480 19456
rect 57428 18148 57480 18154
rect 57428 18090 57480 18096
rect 57440 17338 57468 18090
rect 57428 17332 57480 17338
rect 57428 17274 57480 17280
rect 57520 17128 57572 17134
rect 57520 17070 57572 17076
rect 57532 15706 57560 17070
rect 57520 15700 57572 15706
rect 57520 15642 57572 15648
rect 57624 14618 57652 22066
rect 57796 22034 57848 22040
rect 57900 21554 57928 24142
rect 58084 23322 58112 24142
rect 58176 23866 58204 30670
rect 58254 30631 58310 30640
rect 58268 30598 58296 30631
rect 58256 30592 58308 30598
rect 58256 30534 58308 30540
rect 58532 26580 58584 26586
rect 58532 26522 58584 26528
rect 58256 26376 58308 26382
rect 58256 26318 58308 26324
rect 58268 25906 58296 26318
rect 58256 25900 58308 25906
rect 58256 25842 58308 25848
rect 58440 25152 58492 25158
rect 58440 25094 58492 25100
rect 58452 24818 58480 25094
rect 58440 24812 58492 24818
rect 58440 24754 58492 24760
rect 58256 24608 58308 24614
rect 58254 24576 58256 24585
rect 58308 24576 58310 24585
rect 58254 24511 58310 24520
rect 58164 23860 58216 23866
rect 58164 23802 58216 23808
rect 58164 23724 58216 23730
rect 58164 23666 58216 23672
rect 58072 23316 58124 23322
rect 58072 23258 58124 23264
rect 58176 22778 58204 23666
rect 58256 23112 58308 23118
rect 58256 23054 58308 23060
rect 58164 22772 58216 22778
rect 58164 22714 58216 22720
rect 58072 22228 58124 22234
rect 58072 22170 58124 22176
rect 57980 22160 58032 22166
rect 57980 22102 58032 22108
rect 57888 21548 57940 21554
rect 57888 21490 57940 21496
rect 57900 21146 57928 21490
rect 57888 21140 57940 21146
rect 57888 21082 57940 21088
rect 57704 20800 57756 20806
rect 57704 20742 57756 20748
rect 57716 20534 57744 20742
rect 57704 20528 57756 20534
rect 57704 20470 57756 20476
rect 57716 20058 57744 20470
rect 57704 20052 57756 20058
rect 57704 19994 57756 20000
rect 57796 18284 57848 18290
rect 57796 18226 57848 18232
rect 57808 17882 57836 18226
rect 57796 17876 57848 17882
rect 57796 17818 57848 17824
rect 57888 17536 57940 17542
rect 57888 17478 57940 17484
rect 57900 16454 57928 17478
rect 57888 16448 57940 16454
rect 57888 16390 57940 16396
rect 57900 14822 57928 16390
rect 57888 14816 57940 14822
rect 57888 14758 57940 14764
rect 57612 14612 57664 14618
rect 57612 14554 57664 14560
rect 57624 14074 57652 14554
rect 57900 14414 57928 14758
rect 57888 14408 57940 14414
rect 57888 14350 57940 14356
rect 57796 14272 57848 14278
rect 57796 14214 57848 14220
rect 57612 14068 57664 14074
rect 57612 14010 57664 14016
rect 57336 14000 57388 14006
rect 57336 13942 57388 13948
rect 57428 12640 57480 12646
rect 57428 12582 57480 12588
rect 57336 12096 57388 12102
rect 57336 12038 57388 12044
rect 57244 10056 57296 10062
rect 57244 9998 57296 10004
rect 57152 9920 57204 9926
rect 57152 9862 57204 9868
rect 57164 8498 57192 9862
rect 57256 9761 57284 9998
rect 57242 9752 57298 9761
rect 57242 9687 57298 9696
rect 57348 8906 57376 12038
rect 57440 11558 57468 12582
rect 57428 11552 57480 11558
rect 57428 11494 57480 11500
rect 57520 11008 57572 11014
rect 57520 10950 57572 10956
rect 57532 10713 57560 10950
rect 57518 10704 57574 10713
rect 57518 10639 57574 10648
rect 57428 9988 57480 9994
rect 57428 9930 57480 9936
rect 57336 8900 57388 8906
rect 57336 8842 57388 8848
rect 57152 8492 57204 8498
rect 57152 8434 57204 8440
rect 57164 5914 57192 8434
rect 57348 6866 57376 8842
rect 57440 8090 57468 9930
rect 57624 9926 57652 14010
rect 57808 13802 57836 14214
rect 57796 13796 57848 13802
rect 57796 13738 57848 13744
rect 57900 12918 57928 14350
rect 57992 13326 58020 22102
rect 58084 17252 58112 22170
rect 58268 22094 58296 23054
rect 58268 22066 58388 22094
rect 58164 22024 58216 22030
rect 58164 21966 58216 21972
rect 58176 21690 58204 21966
rect 58164 21684 58216 21690
rect 58164 21626 58216 21632
rect 58360 21554 58388 22066
rect 58348 21548 58400 21554
rect 58348 21490 58400 21496
rect 58360 20330 58388 21490
rect 58348 20324 58400 20330
rect 58348 20266 58400 20272
rect 58348 19168 58400 19174
rect 58348 19110 58400 19116
rect 58360 18766 58388 19110
rect 58348 18760 58400 18766
rect 58348 18702 58400 18708
rect 58256 18624 58308 18630
rect 58256 18566 58308 18572
rect 58268 18465 58296 18566
rect 58254 18456 58310 18465
rect 58254 18391 58310 18400
rect 58084 17224 58204 17252
rect 58072 14272 58124 14278
rect 58072 14214 58124 14220
rect 58084 14074 58112 14214
rect 58072 14068 58124 14074
rect 58072 14010 58124 14016
rect 57980 13320 58032 13326
rect 57980 13262 58032 13268
rect 57888 12912 57940 12918
rect 57888 12854 57940 12860
rect 58072 12436 58124 12442
rect 58072 12378 58124 12384
rect 57888 11552 57940 11558
rect 57888 11494 57940 11500
rect 57900 10962 57928 11494
rect 58084 11354 58112 12378
rect 58072 11348 58124 11354
rect 58072 11290 58124 11296
rect 57900 10934 58020 10962
rect 57992 10470 58020 10934
rect 57980 10464 58032 10470
rect 57980 10406 58032 10412
rect 57992 10062 58020 10406
rect 57980 10056 58032 10062
rect 57980 9998 58032 10004
rect 57612 9920 57664 9926
rect 57612 9862 57664 9868
rect 57428 8084 57480 8090
rect 57428 8026 57480 8032
rect 57992 7750 58020 9998
rect 58084 9654 58112 11290
rect 58072 9648 58124 9654
rect 58072 9590 58124 9596
rect 57980 7744 58032 7750
rect 57980 7686 58032 7692
rect 57888 7200 57940 7206
rect 57888 7142 57940 7148
rect 57900 6905 57928 7142
rect 57886 6896 57942 6905
rect 57336 6860 57388 6866
rect 57886 6831 57942 6840
rect 57336 6802 57388 6808
rect 57520 6384 57572 6390
rect 57520 6326 57572 6332
rect 57152 5908 57204 5914
rect 57152 5850 57204 5856
rect 57532 5166 57560 6326
rect 57992 5302 58020 7686
rect 58072 7404 58124 7410
rect 58072 7346 58124 7352
rect 58084 7002 58112 7346
rect 58072 6996 58124 7002
rect 58072 6938 58124 6944
rect 57980 5296 58032 5302
rect 57980 5238 58032 5244
rect 57520 5160 57572 5166
rect 57520 5102 57572 5108
rect 58176 3194 58204 17224
rect 58256 13184 58308 13190
rect 58256 13126 58308 13132
rect 58268 13025 58296 13126
rect 58254 13016 58310 13025
rect 58254 12951 58310 12960
rect 58256 11552 58308 11558
rect 58256 11494 58308 11500
rect 58268 10810 58296 11494
rect 58256 10804 58308 10810
rect 58256 10746 58308 10752
rect 58360 6390 58388 18702
rect 58452 13977 58480 24754
rect 58438 13968 58494 13977
rect 58438 13903 58494 13912
rect 58440 13320 58492 13326
rect 58440 13262 58492 13268
rect 58452 6458 58480 13262
rect 58544 6798 58572 26522
rect 58532 6792 58584 6798
rect 58532 6734 58584 6740
rect 58440 6452 58492 6458
rect 58440 6394 58492 6400
rect 58348 6384 58400 6390
rect 58348 6326 58400 6332
rect 58544 5914 58572 6734
rect 58532 5908 58584 5914
rect 58532 5850 58584 5856
rect 58164 3188 58216 3194
rect 58164 3130 58216 3136
rect 56980 2746 57100 2774
rect 56980 2650 57008 2746
rect 50896 2644 50948 2650
rect 50896 2586 50948 2592
rect 51632 2644 51684 2650
rect 51632 2586 51684 2592
rect 51908 2644 51960 2650
rect 51908 2586 51960 2592
rect 53472 2644 53524 2650
rect 53472 2586 53524 2592
rect 56968 2644 57020 2650
rect 56968 2586 57020 2592
rect 47124 2576 47176 2582
rect 47124 2518 47176 2524
rect 49240 2576 49292 2582
rect 49240 2518 49292 2524
rect 47032 2440 47084 2446
rect 47032 2382 47084 2388
rect 47136 2106 47164 2518
rect 56980 2446 57008 2586
rect 58176 2446 58204 3130
rect 56968 2440 57020 2446
rect 56968 2382 57020 2388
rect 58164 2440 58216 2446
rect 58164 2382 58216 2388
rect 50160 2304 50212 2310
rect 50160 2246 50212 2252
rect 56048 2304 56100 2310
rect 56048 2246 56100 2252
rect 59912 2304 59964 2310
rect 59912 2246 59964 2252
rect 47124 2100 47176 2106
rect 47124 2042 47176 2048
rect 50172 1306 50200 2246
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50172 1278 50292 1306
rect 50264 800 50292 1278
rect 56060 800 56088 2246
rect 5276 734 5488 762
rect 10966 200 11022 800
rect 16762 200 16818 800
rect 21914 200 21970 800
rect 27710 200 27766 800
rect 33506 200 33562 800
rect 38658 200 38714 800
rect 44454 200 44510 800
rect 50250 200 50306 800
rect 56046 200 56102 800
rect 59924 785 59952 2246
rect 59910 776 59966 785
rect 59910 711 59966 720
<< via2 >>
rect 58254 59880 58310 59936
rect 2778 59200 2834 59256
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 1674 53080 1730 53136
rect 1674 46960 1730 47016
rect 1674 40876 1676 40896
rect 1676 40876 1728 40896
rect 1728 40876 1730 40896
rect 1674 40840 1730 40876
rect 1674 35436 1676 35456
rect 1676 35436 1728 35456
rect 1728 35436 1730 35456
rect 1674 35400 1730 35436
rect 1674 29280 1730 29336
rect 1674 23160 1730 23216
rect 1582 17756 1584 17776
rect 1584 17756 1636 17776
rect 1636 17756 1638 17776
rect 1582 17720 1638 17756
rect 1674 11620 1730 11656
rect 1674 11600 1676 11620
rect 1676 11600 1728 11620
rect 1728 11600 1730 11620
rect 1674 5516 1676 5536
rect 1676 5516 1728 5536
rect 1728 5516 1730 5536
rect 1674 5480 1730 5516
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 27986 57196 27988 57216
rect 27988 57196 28040 57216
rect 28040 57196 28042 57216
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1766 5208 1822 5264
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 27986 57160 28042 57196
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 24582 10784 24638 10840
rect 25410 9016 25466 9072
rect 22650 5616 22706 5672
rect 26606 12044 26608 12064
rect 26608 12044 26660 12064
rect 26660 12044 26662 12064
rect 26606 12008 26662 12044
rect 26330 9832 26386 9888
rect 26606 10376 26662 10432
rect 27526 17584 27582 17640
rect 26882 10956 26884 10976
rect 26884 10956 26936 10976
rect 26936 10956 26938 10976
rect 26882 10920 26938 10956
rect 26054 5480 26110 5536
rect 27434 10104 27490 10160
rect 27618 11076 27674 11112
rect 27618 11056 27620 11076
rect 27620 11056 27672 11076
rect 27672 11056 27674 11076
rect 26790 6840 26846 6896
rect 27066 6976 27122 7032
rect 27618 9696 27674 9752
rect 27618 8916 27620 8936
rect 27620 8916 27672 8936
rect 27672 8916 27674 8936
rect 27618 8880 27674 8916
rect 28354 12164 28410 12200
rect 28354 12144 28356 12164
rect 28356 12144 28408 12164
rect 28408 12144 28410 12164
rect 28262 10920 28318 10976
rect 28722 15272 28778 15328
rect 28722 14068 28778 14104
rect 28722 14048 28724 14068
rect 28724 14048 28776 14068
rect 28776 14048 28778 14068
rect 27894 8744 27950 8800
rect 27618 7404 27674 7440
rect 27618 7384 27620 7404
rect 27620 7384 27672 7404
rect 27672 7384 27674 7404
rect 27342 6160 27398 6216
rect 28538 10412 28540 10432
rect 28540 10412 28592 10432
rect 28592 10412 28594 10432
rect 28078 9832 28134 9888
rect 27986 7384 28042 7440
rect 27986 7284 27988 7304
rect 27988 7284 28040 7304
rect 28040 7284 28042 7304
rect 27986 7248 28042 7284
rect 27618 5344 27674 5400
rect 28538 10376 28594 10412
rect 28446 10260 28502 10296
rect 28446 10240 28448 10260
rect 28448 10240 28500 10260
rect 28500 10240 28502 10260
rect 28262 10104 28318 10160
rect 28262 9052 28264 9072
rect 28264 9052 28316 9072
rect 28316 9052 28318 9072
rect 28262 9016 28318 9052
rect 28354 6996 28410 7032
rect 28354 6976 28356 6996
rect 28356 6976 28408 6996
rect 28408 6976 28410 6996
rect 28906 10920 28962 10976
rect 28906 9152 28962 9208
rect 29274 10532 29330 10568
rect 29274 10512 29276 10532
rect 29276 10512 29328 10532
rect 29328 10512 29330 10532
rect 29182 9560 29238 9616
rect 29090 9016 29146 9072
rect 29090 7928 29146 7984
rect 29642 8916 29644 8936
rect 29644 8916 29696 8936
rect 29696 8916 29698 8936
rect 29642 8880 29698 8916
rect 29458 8336 29514 8392
rect 29182 6840 29238 6896
rect 28722 6024 28778 6080
rect 29274 6024 29330 6080
rect 28446 5480 28502 5536
rect 28538 5072 28594 5128
rect 28906 5480 28962 5536
rect 28722 5344 28778 5400
rect 28630 4936 28686 4992
rect 27986 4020 27988 4040
rect 27988 4020 28040 4040
rect 28040 4020 28042 4040
rect 27986 3984 28042 4020
rect 29458 7656 29514 7712
rect 30286 11736 30342 11792
rect 30194 11192 30250 11248
rect 30378 11328 30434 11384
rect 30286 10804 30342 10840
rect 30286 10784 30288 10804
rect 30288 10784 30340 10804
rect 30340 10784 30342 10804
rect 30102 10512 30158 10568
rect 29918 10104 29974 10160
rect 29826 9580 29882 9616
rect 29826 9560 29828 9580
rect 29828 9560 29880 9580
rect 29880 9560 29882 9580
rect 29826 8880 29882 8936
rect 30010 9152 30066 9208
rect 30010 9036 30066 9072
rect 30010 9016 30012 9036
rect 30012 9016 30064 9036
rect 30064 9016 30066 9036
rect 30286 8608 30342 8664
rect 30286 8372 30288 8392
rect 30288 8372 30340 8392
rect 30340 8372 30342 8392
rect 30286 8336 30342 8372
rect 30010 7928 30066 7984
rect 29826 6432 29882 6488
rect 29918 5616 29974 5672
rect 30102 7384 30158 7440
rect 31574 16632 31630 16688
rect 31022 13776 31078 13832
rect 31022 11600 31078 11656
rect 30930 10512 30986 10568
rect 30930 10104 30986 10160
rect 31206 9988 31262 10024
rect 31206 9968 31208 9988
rect 31208 9968 31260 9988
rect 31260 9968 31262 9988
rect 30930 8744 30986 8800
rect 31574 11600 31630 11656
rect 31850 11192 31906 11248
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 31942 11056 31998 11112
rect 31758 10104 31814 10160
rect 31206 7520 31262 7576
rect 31114 7384 31170 7440
rect 30102 5364 30158 5400
rect 30102 5344 30104 5364
rect 30104 5344 30156 5364
rect 30156 5344 30158 5364
rect 31390 8492 31446 8528
rect 31390 8472 31392 8492
rect 31392 8472 31444 8492
rect 31444 8472 31446 8492
rect 31758 7928 31814 7984
rect 31666 7384 31722 7440
rect 31666 6976 31722 7032
rect 31850 6976 31906 7032
rect 32310 11056 32366 11112
rect 32494 11756 32550 11792
rect 32494 11736 32496 11756
rect 32496 11736 32548 11756
rect 32548 11736 32550 11756
rect 32126 9560 32182 9616
rect 32310 9424 32366 9480
rect 32310 8900 32366 8936
rect 32310 8880 32312 8900
rect 32312 8880 32364 8900
rect 32364 8880 32366 8900
rect 32126 8472 32182 8528
rect 32034 8200 32090 8256
rect 31390 6024 31446 6080
rect 31390 5908 31446 5944
rect 31390 5888 31392 5908
rect 31392 5888 31444 5908
rect 31444 5888 31446 5908
rect 32126 6452 32182 6488
rect 32126 6432 32128 6452
rect 32128 6432 32180 6452
rect 32180 6432 32182 6452
rect 32494 8880 32550 8936
rect 32494 7384 32550 7440
rect 32494 6704 32550 6760
rect 32770 11076 32826 11112
rect 32770 11056 32772 11076
rect 32772 11056 32824 11076
rect 32824 11056 32826 11076
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 33322 12300 33378 12336
rect 33322 12280 33324 12300
rect 33324 12280 33376 12300
rect 33376 12280 33378 12300
rect 33322 10920 33378 10976
rect 32954 9696 33010 9752
rect 33322 9696 33378 9752
rect 33046 9424 33102 9480
rect 32770 8744 32826 8800
rect 32770 8064 32826 8120
rect 32586 6160 32642 6216
rect 33230 7148 33232 7168
rect 33232 7148 33284 7168
rect 33284 7148 33286 7168
rect 33230 7112 33286 7148
rect 33966 12144 34022 12200
rect 33782 11348 33838 11384
rect 33782 11328 33784 11348
rect 33784 11328 33836 11348
rect 33836 11328 33838 11348
rect 33690 9988 33746 10024
rect 33690 9968 33692 9988
rect 33692 9968 33744 9988
rect 33744 9968 33746 9988
rect 34242 10548 34244 10568
rect 34244 10548 34296 10568
rect 34296 10548 34298 10568
rect 34242 10512 34298 10548
rect 34150 10240 34206 10296
rect 34150 9832 34206 9888
rect 34058 9696 34114 9752
rect 33506 6568 33562 6624
rect 34150 7792 34206 7848
rect 33782 6568 33838 6624
rect 33782 5364 33838 5400
rect 33782 5344 33784 5364
rect 33784 5344 33836 5364
rect 33836 5344 33838 5364
rect 33874 4936 33930 4992
rect 34150 6160 34206 6216
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34886 14048 34942 14104
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34978 12688 35034 12744
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 36082 20204 36084 20224
rect 36084 20204 36136 20224
rect 36136 20204 36138 20224
rect 36082 20168 36138 20204
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35622 11056 35678 11112
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34518 8064 34574 8120
rect 35254 8492 35310 8528
rect 35254 8472 35256 8492
rect 35256 8472 35308 8492
rect 35308 8472 35310 8492
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35162 7948 35218 7984
rect 35162 7928 35164 7948
rect 35164 7928 35216 7948
rect 35216 7928 35218 7948
rect 35806 9424 35862 9480
rect 35622 7540 35678 7576
rect 35898 8744 35954 8800
rect 35990 7928 36046 7984
rect 35622 7520 35624 7540
rect 35624 7520 35676 7540
rect 35676 7520 35678 7540
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34334 5072 34390 5128
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35530 7268 35586 7304
rect 35530 7248 35532 7268
rect 35532 7248 35584 7268
rect 35584 7248 35586 7268
rect 35070 5344 35126 5400
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36726 11756 36782 11792
rect 36726 11736 36728 11756
rect 36728 11736 36780 11756
rect 36780 11736 36782 11756
rect 36174 8880 36230 8936
rect 37002 12724 37004 12744
rect 37004 12724 37056 12744
rect 37056 12724 37058 12744
rect 37002 12688 37058 12724
rect 36910 11076 36966 11112
rect 36910 11056 36912 11076
rect 36912 11056 36964 11076
rect 36964 11056 36966 11076
rect 36818 9288 36874 9344
rect 36082 6840 36138 6896
rect 36450 6840 36506 6896
rect 37278 9424 37334 9480
rect 38934 17040 38990 17096
rect 37646 12180 37648 12200
rect 37648 12180 37700 12200
rect 37700 12180 37702 12200
rect 37646 12144 37702 12180
rect 37554 11620 37610 11656
rect 37554 11600 37556 11620
rect 37556 11600 37608 11620
rect 37608 11600 37610 11620
rect 37278 8372 37280 8392
rect 37280 8372 37332 8392
rect 37332 8372 37334 8392
rect 37278 8336 37334 8372
rect 37646 9324 37648 9344
rect 37648 9324 37700 9344
rect 37700 9324 37702 9344
rect 37646 9288 37702 9324
rect 35714 5072 35770 5128
rect 36082 4548 36138 4584
rect 36082 4528 36084 4548
rect 36084 4528 36136 4548
rect 36136 4528 36138 4548
rect 37278 5480 37334 5536
rect 38198 9444 38254 9480
rect 38198 9424 38200 9444
rect 38200 9424 38252 9444
rect 38252 9424 38254 9444
rect 39854 13776 39910 13832
rect 40498 13776 40554 13832
rect 38842 9172 38898 9208
rect 38842 9152 38844 9172
rect 38844 9152 38896 9172
rect 38896 9152 38898 9172
rect 40406 12280 40462 12336
rect 38382 7792 38438 7848
rect 37922 6432 37978 6488
rect 37830 5480 37886 5536
rect 38014 5344 38070 5400
rect 38658 6332 38660 6352
rect 38660 6332 38712 6352
rect 38712 6332 38714 6352
rect 38658 6296 38714 6332
rect 38290 5752 38346 5808
rect 40406 6316 40462 6352
rect 40406 6296 40408 6316
rect 40408 6296 40460 6316
rect 40460 6296 40462 6316
rect 41326 10004 41328 10024
rect 41328 10004 41380 10024
rect 41380 10004 41382 10024
rect 41326 9968 41382 10004
rect 41326 9560 41382 9616
rect 41418 5228 41474 5264
rect 41418 5208 41420 5228
rect 41420 5208 41472 5228
rect 41472 5208 41474 5228
rect 41510 4004 41566 4040
rect 41510 3984 41512 4004
rect 41512 3984 41564 4004
rect 41564 3984 41566 4004
rect 42154 4684 42210 4720
rect 42154 4664 42156 4684
rect 42156 4664 42208 4684
rect 42208 4664 42210 4684
rect 43626 19372 43682 19408
rect 43626 19352 43628 19372
rect 43628 19352 43680 19372
rect 43680 19352 43682 19372
rect 43902 18028 43904 18048
rect 43904 18028 43956 18048
rect 43956 18028 43958 18048
rect 43902 17992 43958 18028
rect 43626 15972 43682 16008
rect 43626 15952 43628 15972
rect 43628 15952 43680 15972
rect 43680 15952 43682 15972
rect 42890 13232 42946 13288
rect 43810 13268 43812 13288
rect 43812 13268 43864 13288
rect 43864 13268 43866 13288
rect 43810 13232 43866 13268
rect 43718 13096 43774 13152
rect 44454 20304 44510 20360
rect 43718 12588 43720 12608
rect 43720 12588 43772 12608
rect 43772 12588 43774 12608
rect 43718 12552 43774 12588
rect 43350 9696 43406 9752
rect 43258 5752 43314 5808
rect 43718 9424 43774 9480
rect 43718 7112 43774 7168
rect 43994 12552 44050 12608
rect 44362 16224 44418 16280
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 44454 15544 44510 15600
rect 44362 13640 44418 13696
rect 43994 10956 43996 10976
rect 43996 10956 44048 10976
rect 44048 10956 44050 10976
rect 43994 10920 44050 10956
rect 44270 11892 44326 11928
rect 44270 11872 44272 11892
rect 44272 11872 44324 11892
rect 44324 11872 44326 11892
rect 44362 9696 44418 9752
rect 43902 6840 43958 6896
rect 44914 15020 44970 15056
rect 44914 15000 44916 15020
rect 44916 15000 44968 15020
rect 44968 15000 44970 15020
rect 45282 17040 45338 17096
rect 45006 13504 45062 13560
rect 45006 12144 45062 12200
rect 46110 22516 46112 22536
rect 46112 22516 46164 22536
rect 46164 22516 46166 22536
rect 46110 22480 46166 22516
rect 45742 17720 45798 17776
rect 45466 17620 45468 17640
rect 45468 17620 45520 17640
rect 45520 17620 45522 17640
rect 45466 17584 45522 17620
rect 45190 15816 45246 15872
rect 45926 16088 45982 16144
rect 46110 16360 46166 16416
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50066 27648 50122 27704
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 45374 15408 45430 15464
rect 45282 15308 45284 15328
rect 45284 15308 45336 15328
rect 45336 15308 45338 15328
rect 45282 15272 45338 15308
rect 45282 14864 45338 14920
rect 45374 13096 45430 13152
rect 45190 11872 45246 11928
rect 44822 9288 44878 9344
rect 46202 15408 46258 15464
rect 45558 14320 45614 14376
rect 46938 21292 46940 21312
rect 46940 21292 46992 21312
rect 46992 21292 46994 21312
rect 46938 21256 46994 21292
rect 45742 13368 45798 13424
rect 45466 12180 45468 12200
rect 45468 12180 45520 12200
rect 45520 12180 45522 12200
rect 45466 12144 45522 12180
rect 45282 9968 45338 10024
rect 45650 11872 45706 11928
rect 45558 11056 45614 11112
rect 45834 12688 45890 12744
rect 46202 13232 46258 13288
rect 46202 12688 46258 12744
rect 46386 12144 46442 12200
rect 45742 10784 45798 10840
rect 44546 7812 44602 7848
rect 44546 7792 44548 7812
rect 44548 7792 44600 7812
rect 44600 7792 44602 7812
rect 45926 10260 45982 10296
rect 45926 10240 45928 10260
rect 45928 10240 45980 10260
rect 45980 10240 45982 10260
rect 45650 8880 45706 8936
rect 45374 8492 45430 8528
rect 45374 8472 45376 8492
rect 45376 8472 45428 8492
rect 45428 8472 45430 8492
rect 45650 8744 45706 8800
rect 44454 4664 44510 4720
rect 45190 4800 45246 4856
rect 45834 9580 45890 9616
rect 45834 9560 45836 9580
rect 45836 9560 45888 9580
rect 45888 9560 45890 9580
rect 46110 11056 46166 11112
rect 46018 8880 46074 8936
rect 46294 9424 46350 9480
rect 46846 15544 46902 15600
rect 46662 14900 46664 14920
rect 46664 14900 46716 14920
rect 46716 14900 46718 14920
rect 46662 14864 46718 14900
rect 46662 14320 46718 14376
rect 46846 15136 46902 15192
rect 48502 24792 48558 24848
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 47214 16244 47270 16280
rect 47214 16224 47216 16244
rect 47216 16224 47268 16244
rect 47268 16224 47270 16244
rect 47398 16632 47454 16688
rect 47306 16088 47362 16144
rect 47582 17584 47638 17640
rect 46662 13776 46718 13832
rect 46754 13096 46810 13152
rect 46570 12280 46626 12336
rect 46294 9016 46350 9072
rect 47030 13096 47086 13152
rect 47398 13640 47454 13696
rect 46846 10104 46902 10160
rect 46018 5616 46074 5672
rect 46386 5072 46442 5128
rect 47214 11872 47270 11928
rect 47030 9052 47032 9072
rect 47032 9052 47084 9072
rect 47084 9052 47086 9072
rect 47030 9016 47086 9052
rect 47398 9288 47454 9344
rect 47306 8880 47362 8936
rect 46754 7248 46810 7304
rect 49146 20884 49148 20904
rect 49148 20884 49200 20904
rect 49200 20884 49202 20904
rect 49146 20848 49202 20884
rect 48318 17060 48374 17096
rect 48318 17040 48320 17060
rect 48320 17040 48372 17060
rect 48372 17040 48374 17060
rect 48502 17076 48504 17096
rect 48504 17076 48556 17096
rect 48556 17076 48558 17096
rect 48502 17040 48558 17076
rect 48318 16224 48374 16280
rect 47950 15816 48006 15872
rect 47858 15544 47914 15600
rect 47766 15136 47822 15192
rect 48042 13524 48098 13560
rect 48042 13504 48044 13524
rect 48044 13504 48096 13524
rect 48096 13504 48098 13524
rect 48502 15816 48558 15872
rect 48410 15680 48466 15736
rect 48502 14728 48558 14784
rect 48502 14320 48558 14376
rect 48226 13640 48282 13696
rect 47858 13096 47914 13152
rect 47582 8880 47638 8936
rect 48502 13524 48558 13560
rect 48502 13504 48504 13524
rect 48504 13504 48556 13524
rect 48556 13504 48558 13524
rect 48778 16652 48834 16688
rect 48778 16632 48780 16652
rect 48780 16632 48832 16652
rect 48832 16632 48834 16652
rect 48778 15816 48834 15872
rect 48962 16224 49018 16280
rect 48778 14728 48834 14784
rect 48962 14320 49018 14376
rect 48594 13232 48650 13288
rect 48318 12416 48374 12472
rect 48410 12280 48466 12336
rect 48226 10956 48228 10976
rect 48228 10956 48280 10976
rect 48280 10956 48282 10976
rect 48226 10920 48282 10956
rect 47674 7828 47676 7848
rect 47676 7828 47728 7848
rect 47728 7828 47730 7848
rect 47674 7792 47730 7828
rect 47674 6296 47730 6352
rect 48318 8472 48374 8528
rect 48318 8200 48374 8256
rect 48594 12180 48596 12200
rect 48596 12180 48648 12200
rect 48648 12180 48650 12200
rect 48594 12144 48650 12180
rect 49054 12552 49110 12608
rect 48962 12300 49018 12336
rect 48962 12280 48964 12300
rect 48964 12280 49016 12300
rect 49016 12280 49018 12300
rect 49238 16360 49294 16416
rect 49238 15428 49294 15464
rect 49238 15408 49240 15428
rect 49240 15408 49292 15428
rect 49292 15408 49294 15428
rect 49330 14884 49386 14920
rect 49330 14864 49332 14884
rect 49332 14864 49384 14884
rect 49384 14864 49386 14884
rect 49514 15408 49570 15464
rect 49330 13776 49386 13832
rect 48778 10104 48834 10160
rect 48594 9968 48650 10024
rect 48502 9424 48558 9480
rect 46570 5208 46626 5264
rect 46662 4664 46718 4720
rect 47030 4936 47086 4992
rect 48318 6840 48374 6896
rect 47674 4936 47730 4992
rect 47398 4820 47454 4856
rect 47398 4800 47400 4820
rect 47400 4800 47452 4820
rect 47452 4800 47454 4820
rect 47582 4392 47638 4448
rect 47950 4392 48006 4448
rect 48686 9288 48742 9344
rect 48962 9152 49018 9208
rect 48870 6976 48926 7032
rect 48502 5092 48558 5128
rect 48502 5072 48504 5092
rect 48504 5072 48556 5092
rect 48556 5072 48558 5092
rect 47030 2644 47086 2680
rect 47030 2624 47032 2644
rect 47032 2624 47084 2644
rect 47084 2624 47086 2644
rect 49422 12844 49478 12880
rect 49422 12824 49424 12844
rect 49424 12824 49476 12844
rect 49476 12824 49478 12844
rect 49606 13676 49608 13696
rect 49608 13676 49660 13696
rect 49660 13676 49662 13696
rect 49606 13640 49662 13676
rect 49698 13388 49754 13424
rect 49698 13368 49700 13388
rect 49700 13368 49752 13388
rect 49752 13368 49754 13388
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50434 17196 50490 17232
rect 50434 17176 50436 17196
rect 50436 17176 50488 17196
rect 50488 17176 50490 17196
rect 50526 17040 50582 17096
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50986 16496 51042 16552
rect 50158 15816 50214 15872
rect 49974 15544 50030 15600
rect 50066 15000 50122 15056
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50250 14864 50306 14920
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 49698 11076 49754 11112
rect 49698 11056 49700 11076
rect 49700 11056 49752 11076
rect 49752 11056 49754 11076
rect 49514 10376 49570 10432
rect 49422 10004 49424 10024
rect 49424 10004 49476 10024
rect 49476 10004 49478 10024
rect 49422 9968 49478 10004
rect 49606 8492 49662 8528
rect 49606 8472 49608 8492
rect 49608 8472 49660 8492
rect 49660 8472 49662 8492
rect 49790 10412 49792 10432
rect 49792 10412 49844 10432
rect 49844 10412 49846 10432
rect 49790 10376 49846 10412
rect 49330 7656 49386 7712
rect 49606 7384 49662 7440
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50342 12552 50398 12608
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50894 14456 50950 14512
rect 51354 16532 51356 16552
rect 51356 16532 51408 16552
rect 51408 16532 51410 16552
rect 51354 16496 51410 16532
rect 51262 16088 51318 16144
rect 50802 12144 50858 12200
rect 50986 12008 51042 12064
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50066 9152 50122 9208
rect 49882 7656 49938 7712
rect 49790 6704 49846 6760
rect 49606 5752 49662 5808
rect 49698 5616 49754 5672
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 51538 15816 51594 15872
rect 51998 19252 52000 19272
rect 52000 19252 52052 19272
rect 52052 19252 52054 19272
rect 51998 19216 52054 19252
rect 51262 12280 51318 12336
rect 51906 14728 51962 14784
rect 53102 17176 53158 17232
rect 52550 15952 52606 16008
rect 52458 15000 52514 15056
rect 50618 8472 50674 8528
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50342 6740 50344 6760
rect 50344 6740 50396 6760
rect 50396 6740 50398 6760
rect 50342 6704 50398 6740
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50342 6316 50398 6352
rect 50342 6296 50344 6316
rect 50344 6296 50396 6316
rect 50396 6296 50398 6316
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 51538 9424 51594 9480
rect 51354 8472 51410 8528
rect 51078 7284 51080 7304
rect 51080 7284 51132 7304
rect 51132 7284 51134 7304
rect 51078 7248 51134 7284
rect 52182 11192 52238 11248
rect 52182 10512 52238 10568
rect 51814 8084 51870 8120
rect 51814 8064 51816 8084
rect 51816 8064 51868 8084
rect 51868 8064 51870 8084
rect 52182 9560 52238 9616
rect 52366 13504 52422 13560
rect 53194 16632 53250 16688
rect 52366 12180 52368 12200
rect 52368 12180 52420 12200
rect 52420 12180 52422 12200
rect 52366 12144 52422 12180
rect 52366 10920 52422 10976
rect 51170 6316 51226 6352
rect 51170 6296 51172 6316
rect 51172 6296 51224 6316
rect 51224 6296 51226 6316
rect 51722 6316 51778 6352
rect 51722 6296 51724 6316
rect 51724 6296 51776 6316
rect 51776 6296 51778 6316
rect 51538 5208 51594 5264
rect 51630 4528 51686 4584
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 54022 17992 54078 18048
rect 53470 14884 53526 14920
rect 53470 14864 53472 14884
rect 53472 14864 53524 14884
rect 53524 14864 53526 14884
rect 53102 13232 53158 13288
rect 52734 11600 52790 11656
rect 52458 9696 52514 9752
rect 52458 9580 52514 9616
rect 52458 9560 52460 9580
rect 52460 9560 52512 9580
rect 52512 9560 52514 9580
rect 53838 15000 53894 15056
rect 54298 16496 54354 16552
rect 53378 12316 53380 12336
rect 53380 12316 53432 12336
rect 53432 12316 53434 12336
rect 53378 12280 53434 12316
rect 53102 11092 53104 11112
rect 53104 11092 53156 11112
rect 53156 11092 53158 11112
rect 53102 11056 53158 11092
rect 52550 9288 52606 9344
rect 52550 8880 52606 8936
rect 53654 12144 53710 12200
rect 53470 9696 53526 9752
rect 53378 6976 53434 7032
rect 53654 9968 53710 10024
rect 53746 9560 53802 9616
rect 54206 12416 54262 12472
rect 55218 15136 55274 15192
rect 55586 15680 55642 15736
rect 55218 14456 55274 14512
rect 54758 12416 54814 12472
rect 54022 10804 54078 10840
rect 54022 10784 54024 10804
rect 54024 10784 54076 10804
rect 54076 10784 54078 10804
rect 54298 10920 54354 10976
rect 54666 10376 54722 10432
rect 54206 8200 54262 8256
rect 54850 6724 54906 6760
rect 54850 6704 54852 6724
rect 54852 6704 54904 6724
rect 54904 6704 54906 6724
rect 55402 12588 55404 12608
rect 55404 12588 55456 12608
rect 55456 12588 55458 12608
rect 55402 12552 55458 12588
rect 55126 10804 55182 10840
rect 55126 10784 55128 10804
rect 55128 10784 55180 10804
rect 55180 10784 55182 10804
rect 55494 12316 55496 12336
rect 55496 12316 55548 12336
rect 55548 12316 55550 12336
rect 55494 12280 55550 12316
rect 55218 7384 55274 7440
rect 56598 13524 56654 13560
rect 56598 13504 56600 13524
rect 56600 13504 56652 13524
rect 56652 13504 56654 13524
rect 56598 10648 56654 10704
rect 56414 8880 56470 8936
rect 58254 54476 58256 54496
rect 58256 54476 58308 54496
rect 58308 54476 58310 54496
rect 58254 54440 58310 54476
rect 58254 48320 58310 48376
rect 58254 42200 58310 42256
rect 58254 36760 58310 36816
rect 58254 30640 58310 30696
rect 58254 24556 58256 24576
rect 58256 24556 58308 24576
rect 58308 24556 58310 24576
rect 58254 24520 58310 24556
rect 57242 9696 57298 9752
rect 57518 10648 57574 10704
rect 58254 18400 58310 18456
rect 57886 6840 57942 6896
rect 58254 12960 58310 13016
rect 58438 13912 58494 13968
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 59910 720 59966 776
<< metal3 >>
rect 58249 59938 58315 59941
rect 59200 59938 59800 59968
rect 58249 59936 59800 59938
rect 58249 59880 58254 59936
rect 58310 59880 59800 59936
rect 58249 59878 59800 59880
rect 58249 59875 58315 59878
rect 59200 59848 59800 59878
rect 200 59258 800 59288
rect 2773 59258 2839 59261
rect 200 59256 2839 59258
rect 200 59200 2778 59256
rect 2834 59200 2839 59256
rect 200 59198 2839 59200
rect 200 59168 800 59198
rect 2773 59195 2839 59198
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 27981 57220 28047 57221
rect 27981 57218 28028 57220
rect 27936 57216 28028 57218
rect 27936 57160 27986 57216
rect 27936 57158 28028 57160
rect 27981 57156 28028 57158
rect 28092 57156 28098 57220
rect 27981 57155 28047 57156
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 58249 54498 58315 54501
rect 59200 54498 59800 54528
rect 58249 54496 59800 54498
rect 58249 54440 58254 54496
rect 58310 54440 59800 54496
rect 58249 54438 59800 54440
rect 58249 54435 58315 54438
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 59200 54408 59800 54438
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 200 53138 800 53168
rect 1669 53138 1735 53141
rect 200 53136 1735 53138
rect 200 53080 1674 53136
rect 1730 53080 1735 53136
rect 200 53078 1735 53080
rect 200 53048 800 53078
rect 1669 53075 1735 53078
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 58249 48378 58315 48381
rect 59200 48378 59800 48408
rect 58249 48376 59800 48378
rect 58249 48320 58254 48376
rect 58310 48320 59800 48376
rect 58249 48318 59800 48320
rect 58249 48315 58315 48318
rect 59200 48288 59800 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 200 47018 800 47048
rect 1669 47018 1735 47021
rect 200 47016 1735 47018
rect 200 46960 1674 47016
rect 1730 46960 1735 47016
rect 200 46958 1735 46960
rect 200 46928 800 46958
rect 1669 46955 1735 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 58249 42258 58315 42261
rect 59200 42258 59800 42288
rect 58249 42256 59800 42258
rect 58249 42200 58254 42256
rect 58310 42200 59800 42256
rect 58249 42198 59800 42200
rect 58249 42195 58315 42198
rect 59200 42168 59800 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 200 40898 800 40928
rect 1669 40898 1735 40901
rect 200 40896 1735 40898
rect 200 40840 1674 40896
rect 1730 40840 1735 40896
rect 200 40838 1735 40840
rect 200 40808 800 40838
rect 1669 40835 1735 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 58249 36818 58315 36821
rect 59200 36818 59800 36848
rect 58249 36816 59800 36818
rect 58249 36760 58254 36816
rect 58310 36760 59800 36816
rect 58249 36758 59800 36760
rect 58249 36755 58315 36758
rect 59200 36728 59800 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 200 35458 800 35488
rect 1669 35458 1735 35461
rect 200 35456 1735 35458
rect 200 35400 1674 35456
rect 1730 35400 1735 35456
rect 200 35398 1735 35400
rect 200 35368 800 35398
rect 1669 35395 1735 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 58249 30698 58315 30701
rect 59200 30698 59800 30728
rect 58249 30696 59800 30698
rect 58249 30640 58254 30696
rect 58310 30640 59800 30696
rect 58249 30638 59800 30640
rect 58249 30635 58315 30638
rect 59200 30608 59800 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 200 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 1669 29338 1735 29341
rect 200 29336 1735 29338
rect 200 29280 1674 29336
rect 1730 29280 1735 29336
rect 200 29278 1735 29280
rect 200 29248 800 29278
rect 1669 29275 1735 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 49918 27644 49924 27708
rect 49988 27706 49994 27708
rect 50061 27706 50127 27709
rect 49988 27704 50127 27706
rect 49988 27648 50066 27704
rect 50122 27648 50127 27704
rect 49988 27646 50127 27648
rect 49988 27644 49994 27646
rect 50061 27643 50127 27646
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 48497 24850 48563 24853
rect 49366 24850 49372 24852
rect 48497 24848 49372 24850
rect 48497 24792 48502 24848
rect 48558 24792 49372 24848
rect 48497 24790 49372 24792
rect 48497 24787 48563 24790
rect 49366 24788 49372 24790
rect 49436 24788 49442 24852
rect 58249 24578 58315 24581
rect 59200 24578 59800 24608
rect 58249 24576 59800 24578
rect 58249 24520 58254 24576
rect 58310 24520 59800 24576
rect 58249 24518 59800 24520
rect 58249 24515 58315 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 59200 24488 59800 24518
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 200 23218 800 23248
rect 1669 23218 1735 23221
rect 200 23216 1735 23218
rect 200 23160 1674 23216
rect 1730 23160 1735 23216
rect 200 23158 1735 23160
rect 200 23128 800 23158
rect 1669 23155 1735 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 46105 22540 46171 22541
rect 46054 22476 46060 22540
rect 46124 22538 46171 22540
rect 46124 22536 46216 22538
rect 46166 22480 46216 22536
rect 46124 22478 46216 22480
rect 46124 22476 46171 22478
rect 46105 22475 46171 22476
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 46933 21314 46999 21317
rect 53414 21314 53420 21316
rect 46933 21312 53420 21314
rect 46933 21256 46938 21312
rect 46994 21256 53420 21312
rect 46933 21254 53420 21256
rect 46933 21251 46999 21254
rect 53414 21252 53420 21254
rect 53484 21252 53490 21316
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 49141 20908 49207 20909
rect 49141 20906 49188 20908
rect 49096 20904 49188 20906
rect 49096 20848 49146 20904
rect 49096 20846 49188 20848
rect 49141 20844 49188 20846
rect 49252 20844 49258 20908
rect 49141 20843 49207 20844
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 44449 20362 44515 20365
rect 44582 20362 44588 20364
rect 44449 20360 44588 20362
rect 44449 20304 44454 20360
rect 44510 20304 44588 20360
rect 44449 20302 44588 20304
rect 44449 20299 44515 20302
rect 44582 20300 44588 20302
rect 44652 20300 44658 20364
rect 36077 20228 36143 20229
rect 36077 20226 36124 20228
rect 36032 20224 36124 20226
rect 36032 20168 36082 20224
rect 36032 20166 36124 20168
rect 36077 20164 36124 20166
rect 36188 20164 36194 20228
rect 36077 20163 36143 20164
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 43621 19412 43687 19413
rect 43621 19410 43668 19412
rect 43576 19408 43668 19410
rect 43576 19352 43626 19408
rect 43576 19350 43668 19352
rect 43621 19348 43668 19350
rect 43732 19348 43738 19412
rect 43621 19347 43687 19348
rect 51993 19274 52059 19277
rect 52310 19274 52316 19276
rect 51993 19272 52316 19274
rect 51993 19216 51998 19272
rect 52054 19216 52316 19272
rect 51993 19214 52316 19216
rect 51993 19211 52059 19214
rect 52310 19212 52316 19214
rect 52380 19212 52386 19276
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 58249 18458 58315 18461
rect 59200 18458 59800 18488
rect 58249 18456 59800 18458
rect 58249 18400 58254 18456
rect 58310 18400 59800 18456
rect 58249 18398 59800 18400
rect 58249 18395 58315 18398
rect 59200 18368 59800 18398
rect 43897 18050 43963 18053
rect 54017 18052 54083 18053
rect 44030 18050 44036 18052
rect 43897 18048 44036 18050
rect 43897 17992 43902 18048
rect 43958 17992 44036 18048
rect 43897 17990 44036 17992
rect 43897 17987 43963 17990
rect 44030 17988 44036 17990
rect 44100 17988 44106 18052
rect 53966 18050 53972 18052
rect 53926 17990 53972 18050
rect 54036 18048 54083 18052
rect 54078 17992 54083 18048
rect 53966 17988 53972 17990
rect 54036 17988 54083 17992
rect 54017 17987 54083 17988
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 200 17778 800 17808
rect 1577 17778 1643 17781
rect 45737 17780 45803 17781
rect 200 17776 1643 17778
rect 200 17720 1582 17776
rect 1638 17720 1643 17776
rect 200 17718 1643 17720
rect 200 17688 800 17718
rect 1577 17715 1643 17718
rect 45686 17716 45692 17780
rect 45756 17778 45803 17780
rect 45756 17776 45848 17778
rect 45798 17720 45848 17776
rect 45756 17718 45848 17720
rect 45756 17716 45803 17718
rect 45737 17715 45803 17716
rect 27521 17644 27587 17645
rect 27470 17580 27476 17644
rect 27540 17642 27587 17644
rect 45461 17642 45527 17645
rect 47577 17642 47643 17645
rect 27540 17640 27632 17642
rect 27582 17584 27632 17640
rect 27540 17582 27632 17584
rect 45461 17640 47643 17642
rect 45461 17584 45466 17640
rect 45522 17584 47582 17640
rect 47638 17584 47643 17640
rect 45461 17582 47643 17584
rect 27540 17580 27587 17582
rect 27521 17579 27587 17580
rect 45461 17579 45527 17582
rect 47577 17579 47643 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 50429 17234 50495 17237
rect 53097 17234 53163 17237
rect 50429 17232 53163 17234
rect 50429 17176 50434 17232
rect 50490 17176 53102 17232
rect 53158 17176 53163 17232
rect 50429 17174 53163 17176
rect 50429 17171 50495 17174
rect 53097 17171 53163 17174
rect 38929 17100 38995 17101
rect 38878 17036 38884 17100
rect 38948 17098 38995 17100
rect 45277 17098 45343 17101
rect 48313 17100 48379 17101
rect 48262 17098 48268 17100
rect 38948 17096 39040 17098
rect 38990 17040 39040 17096
rect 38948 17038 39040 17040
rect 45277 17096 48268 17098
rect 48332 17096 48379 17100
rect 45277 17040 45282 17096
rect 45338 17040 48268 17096
rect 48374 17040 48379 17096
rect 45277 17038 48268 17040
rect 38948 17036 38995 17038
rect 38929 17035 38995 17036
rect 45277 17035 45343 17038
rect 48262 17036 48268 17038
rect 48332 17036 48379 17040
rect 48313 17035 48379 17036
rect 48497 17098 48563 17101
rect 48630 17098 48636 17100
rect 48497 17096 48636 17098
rect 48497 17040 48502 17096
rect 48558 17040 48636 17096
rect 48497 17038 48636 17040
rect 48497 17035 48563 17038
rect 48630 17036 48636 17038
rect 48700 17098 48706 17100
rect 50521 17098 50587 17101
rect 48700 17096 50587 17098
rect 48700 17040 50526 17096
rect 50582 17040 50587 17096
rect 48700 17038 50587 17040
rect 48700 17036 48706 17038
rect 50521 17035 50587 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 31569 16692 31635 16693
rect 31518 16628 31524 16692
rect 31588 16690 31635 16692
rect 47393 16690 47459 16693
rect 48773 16690 48839 16693
rect 31588 16688 31680 16690
rect 31630 16632 31680 16688
rect 31588 16630 31680 16632
rect 47393 16688 48839 16690
rect 47393 16632 47398 16688
rect 47454 16632 48778 16688
rect 48834 16632 48839 16688
rect 47393 16630 48839 16632
rect 31588 16628 31635 16630
rect 31569 16627 31635 16628
rect 47393 16627 47459 16630
rect 48773 16627 48839 16630
rect 53189 16690 53255 16693
rect 53782 16690 53788 16692
rect 53189 16688 53788 16690
rect 53189 16632 53194 16688
rect 53250 16632 53788 16688
rect 53189 16630 53788 16632
rect 53189 16627 53255 16630
rect 53782 16628 53788 16630
rect 53852 16628 53858 16692
rect 49182 16492 49188 16556
rect 49252 16554 49258 16556
rect 50981 16554 51047 16557
rect 49252 16552 51047 16554
rect 49252 16496 50986 16552
rect 51042 16496 51047 16552
rect 49252 16494 51047 16496
rect 49252 16492 49258 16494
rect 50981 16491 51047 16494
rect 51349 16554 51415 16557
rect 54293 16554 54359 16557
rect 51349 16552 54359 16554
rect 51349 16496 51354 16552
rect 51410 16496 54298 16552
rect 54354 16496 54359 16552
rect 51349 16494 54359 16496
rect 51349 16491 51415 16494
rect 54293 16491 54359 16494
rect 46105 16418 46171 16421
rect 49233 16418 49299 16421
rect 46105 16416 49299 16418
rect 46105 16360 46110 16416
rect 46166 16360 49238 16416
rect 49294 16360 49299 16416
rect 46105 16358 49299 16360
rect 46105 16355 46171 16358
rect 49233 16355 49299 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 44357 16282 44423 16285
rect 47209 16282 47275 16285
rect 44357 16280 47275 16282
rect 44357 16224 44362 16280
rect 44418 16224 47214 16280
rect 47270 16224 47275 16280
rect 44357 16222 47275 16224
rect 44357 16219 44423 16222
rect 47209 16219 47275 16222
rect 48313 16282 48379 16285
rect 48957 16282 49023 16285
rect 48313 16280 49023 16282
rect 48313 16224 48318 16280
rect 48374 16224 48962 16280
rect 49018 16224 49023 16280
rect 48313 16222 49023 16224
rect 48313 16219 48379 16222
rect 48957 16219 49023 16222
rect 45921 16146 45987 16149
rect 47301 16146 47367 16149
rect 51257 16146 51323 16149
rect 45921 16144 51323 16146
rect 45921 16088 45926 16144
rect 45982 16088 47306 16144
rect 47362 16088 51262 16144
rect 51318 16088 51323 16144
rect 45921 16086 51323 16088
rect 45921 16083 45987 16086
rect 47301 16083 47367 16086
rect 51257 16083 51323 16086
rect 43621 16010 43687 16013
rect 52545 16010 52611 16013
rect 43621 16008 52611 16010
rect 43621 15952 43626 16008
rect 43682 15952 52550 16008
rect 52606 15952 52611 16008
rect 43621 15950 52611 15952
rect 43621 15947 43687 15950
rect 52545 15947 52611 15950
rect 45185 15874 45251 15877
rect 47945 15874 48011 15877
rect 45185 15872 48011 15874
rect 45185 15816 45190 15872
rect 45246 15816 47950 15872
rect 48006 15816 48011 15872
rect 45185 15814 48011 15816
rect 45185 15811 45251 15814
rect 47945 15811 48011 15814
rect 48497 15874 48563 15877
rect 48773 15874 48839 15877
rect 48497 15872 48839 15874
rect 48497 15816 48502 15872
rect 48558 15816 48778 15872
rect 48834 15816 48839 15872
rect 48497 15814 48839 15816
rect 48497 15811 48563 15814
rect 48773 15811 48839 15814
rect 50153 15874 50219 15877
rect 51533 15874 51599 15877
rect 50153 15872 51599 15874
rect 50153 15816 50158 15872
rect 50214 15816 51538 15872
rect 51594 15816 51599 15872
rect 50153 15814 51599 15816
rect 50153 15811 50219 15814
rect 51533 15811 51599 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 48405 15738 48471 15741
rect 55581 15738 55647 15741
rect 48405 15736 55647 15738
rect 48405 15680 48410 15736
rect 48466 15680 55586 15736
rect 55642 15680 55647 15736
rect 48405 15678 55647 15680
rect 48405 15675 48471 15678
rect 55581 15675 55647 15678
rect 44449 15602 44515 15605
rect 46841 15602 46907 15605
rect 44449 15600 46907 15602
rect 44449 15544 44454 15600
rect 44510 15544 46846 15600
rect 46902 15544 46907 15600
rect 44449 15542 46907 15544
rect 44449 15539 44515 15542
rect 46841 15539 46907 15542
rect 47853 15602 47919 15605
rect 49969 15602 50035 15605
rect 47853 15600 50035 15602
rect 47853 15544 47858 15600
rect 47914 15544 49974 15600
rect 50030 15544 50035 15600
rect 47853 15542 50035 15544
rect 47853 15539 47919 15542
rect 49969 15539 50035 15542
rect 45369 15468 45435 15469
rect 45318 15404 45324 15468
rect 45388 15466 45435 15468
rect 46197 15466 46263 15469
rect 49233 15468 49299 15469
rect 45388 15464 46263 15466
rect 45430 15408 46202 15464
rect 46258 15408 46263 15464
rect 45388 15406 46263 15408
rect 45388 15404 45435 15406
rect 45369 15403 45435 15404
rect 46197 15403 46263 15406
rect 49182 15404 49188 15468
rect 49252 15466 49299 15468
rect 49509 15466 49575 15469
rect 49252 15464 49575 15466
rect 49294 15408 49514 15464
rect 49570 15408 49575 15464
rect 49252 15406 49575 15408
rect 49252 15404 49299 15406
rect 49233 15403 49299 15404
rect 49509 15403 49575 15406
rect 28717 15330 28783 15333
rect 30230 15330 30236 15332
rect 28717 15328 30236 15330
rect 28717 15272 28722 15328
rect 28778 15272 30236 15328
rect 28717 15270 30236 15272
rect 28717 15267 28783 15270
rect 30230 15268 30236 15270
rect 30300 15268 30306 15332
rect 45277 15330 45343 15333
rect 45502 15330 45508 15332
rect 45277 15328 45508 15330
rect 45277 15272 45282 15328
rect 45338 15272 45508 15328
rect 45277 15270 45508 15272
rect 45277 15267 45343 15270
rect 45502 15268 45508 15270
rect 45572 15268 45578 15332
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 46841 15194 46907 15197
rect 47761 15194 47827 15197
rect 46841 15192 47827 15194
rect 46841 15136 46846 15192
rect 46902 15136 47766 15192
rect 47822 15136 47827 15192
rect 46841 15134 47827 15136
rect 46841 15131 46907 15134
rect 47761 15131 47827 15134
rect 53414 15132 53420 15196
rect 53484 15194 53490 15196
rect 55213 15194 55279 15197
rect 53484 15192 55279 15194
rect 53484 15136 55218 15192
rect 55274 15136 55279 15192
rect 53484 15134 55279 15136
rect 53484 15132 53490 15134
rect 55213 15131 55279 15134
rect 44909 15058 44975 15061
rect 50061 15058 50127 15061
rect 52453 15058 52519 15061
rect 53833 15058 53899 15061
rect 44909 15056 53899 15058
rect 44909 15000 44914 15056
rect 44970 15000 50066 15056
rect 50122 15000 52458 15056
rect 52514 15000 53838 15056
rect 53894 15000 53899 15056
rect 44909 14998 53899 15000
rect 44909 14995 44975 14998
rect 50061 14995 50127 14998
rect 52453 14995 52519 14998
rect 53833 14995 53899 14998
rect 45277 14922 45343 14925
rect 46657 14922 46723 14925
rect 49325 14924 49391 14925
rect 49325 14922 49372 14924
rect 45277 14920 46723 14922
rect 45277 14864 45282 14920
rect 45338 14864 46662 14920
rect 46718 14864 46723 14920
rect 45277 14862 46723 14864
rect 49280 14920 49372 14922
rect 49280 14864 49330 14920
rect 49280 14862 49372 14864
rect 45277 14859 45343 14862
rect 46657 14859 46723 14862
rect 49325 14860 49372 14862
rect 49436 14860 49442 14924
rect 50245 14922 50311 14925
rect 53465 14922 53531 14925
rect 50245 14920 53531 14922
rect 50245 14864 50250 14920
rect 50306 14864 53470 14920
rect 53526 14864 53531 14920
rect 50245 14862 53531 14864
rect 49325 14859 49391 14860
rect 50245 14859 50311 14862
rect 53465 14859 53531 14862
rect 48497 14786 48563 14789
rect 48630 14786 48636 14788
rect 48497 14784 48636 14786
rect 48497 14728 48502 14784
rect 48558 14728 48636 14784
rect 48497 14726 48636 14728
rect 48497 14723 48563 14726
rect 48630 14724 48636 14726
rect 48700 14724 48706 14788
rect 48773 14786 48839 14789
rect 51901 14786 51967 14789
rect 48773 14784 51967 14786
rect 48773 14728 48778 14784
rect 48834 14728 51906 14784
rect 51962 14728 51967 14784
rect 48773 14726 51967 14728
rect 48773 14723 48839 14726
rect 51901 14723 51967 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 50889 14514 50955 14517
rect 55213 14514 55279 14517
rect 50889 14512 55279 14514
rect 50889 14456 50894 14512
rect 50950 14456 55218 14512
rect 55274 14456 55279 14512
rect 50889 14454 55279 14456
rect 50889 14451 50955 14454
rect 55213 14451 55279 14454
rect 45553 14378 45619 14381
rect 46657 14378 46723 14381
rect 45553 14376 46723 14378
rect 45553 14320 45558 14376
rect 45614 14320 46662 14376
rect 46718 14320 46723 14376
rect 45553 14318 46723 14320
rect 45553 14315 45619 14318
rect 46657 14315 46723 14318
rect 48497 14378 48563 14381
rect 48957 14378 49023 14381
rect 48497 14376 49023 14378
rect 48497 14320 48502 14376
rect 48558 14320 48962 14376
rect 49018 14320 49023 14376
rect 48497 14318 49023 14320
rect 48497 14315 48563 14318
rect 48957 14315 49023 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 28717 14106 28783 14109
rect 34881 14106 34947 14109
rect 28717 14104 34947 14106
rect 28717 14048 28722 14104
rect 28778 14048 34886 14104
rect 34942 14048 34947 14104
rect 28717 14046 34947 14048
rect 28717 14043 28783 14046
rect 34881 14043 34947 14046
rect 58433 13970 58499 13973
rect 41370 13968 58499 13970
rect 41370 13912 58438 13968
rect 58494 13912 58499 13968
rect 41370 13910 58499 13912
rect 31017 13834 31083 13837
rect 39849 13836 39915 13837
rect 31150 13834 31156 13836
rect 31017 13832 31156 13834
rect 31017 13776 31022 13832
rect 31078 13776 31156 13832
rect 31017 13774 31156 13776
rect 31017 13771 31083 13774
rect 31150 13772 31156 13774
rect 31220 13772 31226 13836
rect 39798 13772 39804 13836
rect 39868 13834 39915 13836
rect 40493 13834 40559 13837
rect 41370 13834 41430 13910
rect 58433 13907 58499 13910
rect 39868 13832 39960 13834
rect 39910 13776 39960 13832
rect 39868 13774 39960 13776
rect 40493 13832 41430 13834
rect 40493 13776 40498 13832
rect 40554 13776 41430 13832
rect 40493 13774 41430 13776
rect 46657 13834 46723 13837
rect 49325 13834 49391 13837
rect 46657 13832 49391 13834
rect 46657 13776 46662 13832
rect 46718 13776 49330 13832
rect 49386 13776 49391 13832
rect 46657 13774 49391 13776
rect 39868 13772 39915 13774
rect 39849 13771 39915 13772
rect 40493 13771 40559 13774
rect 46657 13771 46723 13774
rect 49325 13771 49391 13774
rect 44357 13698 44423 13701
rect 47393 13698 47459 13701
rect 48221 13698 48287 13701
rect 44357 13696 48287 13698
rect 44357 13640 44362 13696
rect 44418 13640 47398 13696
rect 47454 13640 48226 13696
rect 48282 13640 48287 13696
rect 44357 13638 48287 13640
rect 44357 13635 44423 13638
rect 47393 13635 47459 13638
rect 48221 13635 48287 13638
rect 49366 13636 49372 13700
rect 49436 13698 49442 13700
rect 49601 13698 49667 13701
rect 49436 13696 49667 13698
rect 49436 13640 49606 13696
rect 49662 13640 49667 13696
rect 49436 13638 49667 13640
rect 49436 13636 49442 13638
rect 49601 13635 49667 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 45001 13562 45067 13565
rect 48037 13562 48103 13565
rect 48497 13564 48563 13565
rect 48446 13562 48452 13564
rect 45001 13560 48103 13562
rect 45001 13504 45006 13560
rect 45062 13504 48042 13560
rect 48098 13504 48103 13560
rect 45001 13502 48103 13504
rect 48406 13502 48452 13562
rect 48516 13560 48563 13564
rect 48558 13504 48563 13560
rect 45001 13499 45067 13502
rect 48037 13499 48103 13502
rect 48446 13500 48452 13502
rect 48516 13500 48563 13504
rect 48497 13499 48563 13500
rect 52361 13562 52427 13565
rect 56593 13562 56659 13565
rect 52361 13560 56659 13562
rect 52361 13504 52366 13560
rect 52422 13504 56598 13560
rect 56654 13504 56659 13560
rect 52361 13502 56659 13504
rect 52361 13499 52427 13502
rect 56593 13499 56659 13502
rect 45737 13426 45803 13429
rect 49693 13426 49759 13429
rect 45737 13424 49759 13426
rect 45737 13368 45742 13424
rect 45798 13368 49698 13424
rect 49754 13368 49759 13424
rect 45737 13366 49759 13368
rect 45737 13363 45803 13366
rect 49693 13363 49759 13366
rect 42885 13290 42951 13293
rect 43805 13290 43871 13293
rect 46197 13290 46263 13293
rect 42885 13288 46263 13290
rect 42885 13232 42890 13288
rect 42946 13232 43810 13288
rect 43866 13232 46202 13288
rect 46258 13232 46263 13288
rect 42885 13230 46263 13232
rect 42885 13227 42951 13230
rect 43805 13227 43871 13230
rect 46197 13227 46263 13230
rect 48589 13292 48655 13293
rect 48589 13288 48636 13292
rect 48700 13290 48706 13292
rect 53097 13290 53163 13293
rect 48700 13288 53163 13290
rect 48589 13232 48594 13288
rect 48700 13232 53102 13288
rect 53158 13232 53163 13288
rect 48589 13228 48636 13232
rect 48700 13230 53163 13232
rect 48700 13228 48706 13230
rect 48589 13227 48655 13228
rect 53097 13227 53163 13230
rect 43713 13154 43779 13157
rect 45369 13154 45435 13157
rect 46749 13154 46815 13157
rect 43713 13152 43914 13154
rect 43713 13096 43718 13152
rect 43774 13096 43914 13152
rect 43713 13094 43914 13096
rect 43713 13091 43779 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 34973 12746 35039 12749
rect 36997 12746 37063 12749
rect 34973 12744 37063 12746
rect 34973 12688 34978 12744
rect 35034 12688 37002 12744
rect 37058 12688 37063 12744
rect 34973 12686 37063 12688
rect 34973 12683 35039 12686
rect 36997 12683 37063 12686
rect 43713 12610 43779 12613
rect 43854 12610 43914 13094
rect 45369 13152 46815 13154
rect 45369 13096 45374 13152
rect 45430 13096 46754 13152
rect 46810 13096 46815 13152
rect 45369 13094 46815 13096
rect 45369 13091 45435 13094
rect 46749 13091 46815 13094
rect 47025 13154 47091 13157
rect 47342 13154 47348 13156
rect 47025 13152 47348 13154
rect 47025 13096 47030 13152
rect 47086 13096 47348 13152
rect 47025 13094 47348 13096
rect 47025 13091 47091 13094
rect 47342 13092 47348 13094
rect 47412 13154 47418 13156
rect 47853 13154 47919 13157
rect 47412 13152 47919 13154
rect 47412 13096 47858 13152
rect 47914 13096 47919 13152
rect 47412 13094 47919 13096
rect 47412 13092 47418 13094
rect 47853 13091 47919 13094
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 58249 13018 58315 13021
rect 59200 13018 59800 13048
rect 58249 13016 59800 13018
rect 58249 12960 58254 13016
rect 58310 12960 59800 13016
rect 58249 12958 59800 12960
rect 58249 12955 58315 12958
rect 59200 12928 59800 12958
rect 45502 12820 45508 12884
rect 45572 12882 45578 12884
rect 49417 12882 49483 12885
rect 50838 12882 50844 12884
rect 45572 12880 50844 12882
rect 45572 12824 49422 12880
rect 49478 12824 50844 12880
rect 45572 12822 50844 12824
rect 45572 12820 45578 12822
rect 49417 12819 49483 12822
rect 50838 12820 50844 12822
rect 50908 12820 50914 12884
rect 45829 12746 45895 12749
rect 46197 12746 46263 12749
rect 45829 12744 46263 12746
rect 45829 12688 45834 12744
rect 45890 12688 46202 12744
rect 46258 12688 46263 12744
rect 45829 12686 46263 12688
rect 45829 12683 45895 12686
rect 46197 12683 46263 12686
rect 43989 12610 44055 12613
rect 49049 12610 49115 12613
rect 49182 12610 49188 12612
rect 43713 12608 49188 12610
rect 43713 12552 43718 12608
rect 43774 12552 43994 12608
rect 44050 12552 49054 12608
rect 49110 12552 49188 12608
rect 43713 12550 49188 12552
rect 43713 12547 43779 12550
rect 43989 12547 44055 12550
rect 49049 12547 49115 12550
rect 49182 12548 49188 12550
rect 49252 12548 49258 12612
rect 50337 12610 50403 12613
rect 55397 12610 55463 12613
rect 50337 12608 55463 12610
rect 50337 12552 50342 12608
rect 50398 12552 55402 12608
rect 55458 12552 55463 12608
rect 50337 12550 55463 12552
rect 50337 12547 50403 12550
rect 55397 12547 55463 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 48313 12474 48379 12477
rect 54201 12474 54267 12477
rect 54753 12474 54819 12477
rect 48313 12472 54819 12474
rect 48313 12416 48318 12472
rect 48374 12416 54206 12472
rect 54262 12416 54758 12472
rect 54814 12416 54819 12472
rect 48313 12414 54819 12416
rect 48313 12411 48379 12414
rect 54201 12411 54267 12414
rect 54753 12411 54819 12414
rect 33317 12338 33383 12341
rect 40401 12338 40467 12341
rect 46565 12338 46631 12341
rect 33317 12336 40467 12338
rect 33317 12280 33322 12336
rect 33378 12280 40406 12336
rect 40462 12280 40467 12336
rect 33317 12278 40467 12280
rect 33317 12275 33383 12278
rect 40401 12275 40467 12278
rect 46430 12336 46631 12338
rect 46430 12280 46570 12336
rect 46626 12280 46631 12336
rect 46430 12278 46631 12280
rect 46430 12205 46490 12278
rect 46565 12275 46631 12278
rect 48405 12338 48471 12341
rect 48957 12338 49023 12341
rect 51257 12338 51323 12341
rect 48405 12336 51323 12338
rect 48405 12280 48410 12336
rect 48466 12280 48962 12336
rect 49018 12280 51262 12336
rect 51318 12280 51323 12336
rect 48405 12278 51323 12280
rect 48405 12275 48471 12278
rect 48957 12275 49023 12278
rect 51257 12275 51323 12278
rect 52310 12276 52316 12340
rect 52380 12338 52386 12340
rect 53373 12338 53439 12341
rect 52380 12336 53439 12338
rect 52380 12280 53378 12336
rect 53434 12280 53439 12336
rect 52380 12278 53439 12280
rect 52380 12276 52386 12278
rect 53373 12275 53439 12278
rect 53782 12276 53788 12340
rect 53852 12338 53858 12340
rect 55489 12338 55555 12341
rect 53852 12336 55555 12338
rect 53852 12280 55494 12336
rect 55550 12280 55555 12336
rect 53852 12278 55555 12280
rect 53852 12276 53858 12278
rect 55489 12275 55555 12278
rect 28349 12202 28415 12205
rect 29862 12202 29868 12204
rect 28349 12200 29868 12202
rect 28349 12144 28354 12200
rect 28410 12144 29868 12200
rect 28349 12142 29868 12144
rect 28349 12139 28415 12142
rect 29862 12140 29868 12142
rect 29932 12202 29938 12204
rect 33961 12202 34027 12205
rect 37641 12204 37707 12205
rect 37590 12202 37596 12204
rect 29932 12200 34027 12202
rect 29932 12144 33966 12200
rect 34022 12144 34027 12200
rect 29932 12142 34027 12144
rect 37550 12142 37596 12202
rect 37660 12200 37707 12204
rect 37702 12144 37707 12200
rect 29932 12140 29938 12142
rect 33961 12139 34027 12142
rect 37590 12140 37596 12142
rect 37660 12140 37707 12144
rect 37641 12139 37707 12140
rect 45001 12202 45067 12205
rect 45461 12202 45527 12205
rect 45001 12200 45527 12202
rect 45001 12144 45006 12200
rect 45062 12144 45466 12200
rect 45522 12144 45527 12200
rect 45001 12142 45527 12144
rect 45001 12139 45067 12142
rect 45461 12139 45527 12142
rect 46381 12200 46490 12205
rect 46381 12144 46386 12200
rect 46442 12144 46490 12200
rect 46381 12142 46490 12144
rect 46381 12139 46447 12142
rect 48262 12140 48268 12204
rect 48332 12202 48338 12204
rect 48589 12202 48655 12205
rect 48332 12200 48655 12202
rect 48332 12144 48594 12200
rect 48650 12144 48655 12200
rect 48332 12142 48655 12144
rect 48332 12140 48338 12142
rect 48589 12139 48655 12142
rect 50797 12202 50863 12205
rect 52361 12202 52427 12205
rect 53649 12202 53715 12205
rect 50797 12200 50906 12202
rect 50797 12144 50802 12200
rect 50858 12144 50906 12200
rect 50797 12139 50906 12144
rect 52361 12200 53715 12202
rect 52361 12144 52366 12200
rect 52422 12144 53654 12200
rect 53710 12144 53715 12200
rect 52361 12142 53715 12144
rect 52361 12139 52427 12142
rect 53649 12139 53715 12142
rect 26601 12066 26667 12069
rect 26734 12066 26740 12068
rect 26601 12064 26740 12066
rect 26601 12008 26606 12064
rect 26662 12008 26740 12064
rect 26601 12006 26740 12008
rect 26601 12003 26667 12006
rect 26734 12004 26740 12006
rect 26804 12004 26810 12068
rect 50846 12066 50906 12139
rect 50981 12066 51047 12069
rect 50846 12064 51047 12066
rect 50846 12008 50986 12064
rect 51042 12008 51047 12064
rect 50846 12006 51047 12008
rect 50981 12003 51047 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 44030 11868 44036 11932
rect 44100 11930 44106 11932
rect 44265 11930 44331 11933
rect 44100 11928 44331 11930
rect 44100 11872 44270 11928
rect 44326 11872 44331 11928
rect 44100 11870 44331 11872
rect 44100 11868 44106 11870
rect 44265 11867 44331 11870
rect 45185 11930 45251 11933
rect 45645 11930 45711 11933
rect 47209 11930 47275 11933
rect 45185 11928 47275 11930
rect 45185 11872 45190 11928
rect 45246 11872 45650 11928
rect 45706 11872 47214 11928
rect 47270 11872 47275 11928
rect 45185 11870 47275 11872
rect 45185 11867 45251 11870
rect 45645 11867 45711 11870
rect 47209 11867 47275 11870
rect 30281 11794 30347 11797
rect 32489 11794 32555 11797
rect 36721 11794 36787 11797
rect 30281 11792 36787 11794
rect 30281 11736 30286 11792
rect 30342 11736 32494 11792
rect 32550 11736 36726 11792
rect 36782 11736 36787 11792
rect 30281 11734 36787 11736
rect 30281 11731 30347 11734
rect 32489 11731 32555 11734
rect 36721 11731 36787 11734
rect 200 11658 800 11688
rect 1669 11658 1735 11661
rect 200 11656 1735 11658
rect 200 11600 1674 11656
rect 1730 11600 1735 11656
rect 200 11598 1735 11600
rect 200 11568 800 11598
rect 1669 11595 1735 11598
rect 31017 11658 31083 11661
rect 31569 11658 31635 11661
rect 37549 11658 37615 11661
rect 52729 11658 52795 11661
rect 31017 11656 37615 11658
rect 31017 11600 31022 11656
rect 31078 11600 31574 11656
rect 31630 11600 37554 11656
rect 37610 11600 37615 11656
rect 31017 11598 37615 11600
rect 31017 11595 31083 11598
rect 31569 11595 31635 11598
rect 37549 11595 37615 11598
rect 52318 11656 52795 11658
rect 52318 11600 52734 11656
rect 52790 11600 52795 11656
rect 52318 11598 52795 11600
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 30373 11386 30439 11389
rect 33777 11386 33843 11389
rect 30373 11384 33843 11386
rect 30373 11328 30378 11384
rect 30434 11328 33782 11384
rect 33838 11328 33843 11384
rect 30373 11326 33843 11328
rect 30373 11323 30439 11326
rect 33777 11323 33843 11326
rect 30189 11250 30255 11253
rect 31845 11250 31911 11253
rect 30189 11248 31911 11250
rect 30189 11192 30194 11248
rect 30250 11192 31850 11248
rect 31906 11192 31911 11248
rect 30189 11190 31911 11192
rect 30189 11187 30255 11190
rect 31845 11187 31911 11190
rect 52177 11250 52243 11253
rect 52318 11250 52378 11598
rect 52729 11595 52795 11598
rect 52177 11248 52378 11250
rect 52177 11192 52182 11248
rect 52238 11192 52378 11248
rect 52177 11190 52378 11192
rect 52177 11187 52243 11190
rect 27613 11114 27679 11117
rect 27838 11114 27844 11116
rect 27613 11112 27844 11114
rect 27613 11056 27618 11112
rect 27674 11056 27844 11112
rect 27613 11054 27844 11056
rect 27613 11051 27679 11054
rect 27838 11052 27844 11054
rect 27908 11052 27914 11116
rect 31937 11114 32003 11117
rect 32305 11114 32371 11117
rect 31937 11112 32371 11114
rect 31937 11056 31942 11112
rect 31998 11056 32310 11112
rect 32366 11056 32371 11112
rect 31937 11054 32371 11056
rect 31937 11051 32003 11054
rect 32305 11051 32371 11054
rect 32765 11114 32831 11117
rect 35617 11114 35683 11117
rect 32765 11112 35683 11114
rect 32765 11056 32770 11112
rect 32826 11056 35622 11112
rect 35678 11056 35683 11112
rect 32765 11054 35683 11056
rect 32765 11051 32831 11054
rect 35617 11051 35683 11054
rect 35934 11052 35940 11116
rect 36004 11114 36010 11116
rect 36905 11114 36971 11117
rect 36004 11112 36971 11114
rect 36004 11056 36910 11112
rect 36966 11056 36971 11112
rect 36004 11054 36971 11056
rect 36004 11052 36010 11054
rect 36905 11051 36971 11054
rect 45553 11114 45619 11117
rect 46105 11114 46171 11117
rect 45553 11112 46171 11114
rect 45553 11056 45558 11112
rect 45614 11056 46110 11112
rect 46166 11056 46171 11112
rect 45553 11054 46171 11056
rect 45553 11051 45619 11054
rect 46105 11051 46171 11054
rect 49693 11114 49759 11117
rect 53097 11114 53163 11117
rect 49693 11112 53163 11114
rect 49693 11056 49698 11112
rect 49754 11056 53102 11112
rect 53158 11056 53163 11112
rect 49693 11054 53163 11056
rect 49693 11051 49759 11054
rect 53097 11051 53163 11054
rect 26877 10978 26943 10981
rect 28257 10978 28323 10981
rect 28901 10978 28967 10981
rect 33317 10978 33383 10981
rect 26877 10976 28967 10978
rect 26877 10920 26882 10976
rect 26938 10920 28262 10976
rect 28318 10920 28906 10976
rect 28962 10920 28967 10976
rect 26877 10918 28967 10920
rect 26877 10915 26943 10918
rect 28257 10915 28323 10918
rect 28901 10915 28967 10918
rect 31710 10976 33383 10978
rect 31710 10920 33322 10976
rect 33378 10920 33383 10976
rect 31710 10918 33383 10920
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 24577 10842 24643 10845
rect 30281 10842 30347 10845
rect 31710 10842 31770 10918
rect 33317 10915 33383 10918
rect 43989 10978 44055 10981
rect 48221 10978 48287 10981
rect 43989 10976 48287 10978
rect 43989 10920 43994 10976
rect 44050 10920 48226 10976
rect 48282 10920 48287 10976
rect 43989 10918 48287 10920
rect 43989 10915 44055 10918
rect 48221 10915 48287 10918
rect 52361 10978 52427 10981
rect 54293 10978 54359 10981
rect 52361 10976 54359 10978
rect 52361 10920 52366 10976
rect 52422 10920 54298 10976
rect 54354 10920 54359 10976
rect 52361 10918 54359 10920
rect 52361 10915 52427 10918
rect 54293 10915 54359 10918
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 24577 10840 31770 10842
rect 24577 10784 24582 10840
rect 24638 10784 30286 10840
rect 30342 10784 31770 10840
rect 24577 10782 31770 10784
rect 24577 10779 24643 10782
rect 30281 10779 30347 10782
rect 45318 10780 45324 10844
rect 45388 10842 45394 10844
rect 45737 10842 45803 10845
rect 54017 10844 54083 10845
rect 55121 10844 55187 10845
rect 45388 10840 45803 10842
rect 45388 10784 45742 10840
rect 45798 10784 45803 10840
rect 45388 10782 45803 10784
rect 45388 10780 45394 10782
rect 45737 10779 45803 10782
rect 53966 10780 53972 10844
rect 54036 10842 54083 10844
rect 55070 10842 55076 10844
rect 54036 10840 54128 10842
rect 54078 10784 54128 10840
rect 54036 10782 54128 10784
rect 55030 10782 55076 10842
rect 55140 10840 55187 10844
rect 55182 10784 55187 10840
rect 54036 10780 54083 10782
rect 55070 10780 55076 10782
rect 55140 10780 55187 10784
rect 54017 10779 54083 10780
rect 55121 10779 55187 10780
rect 56593 10706 56659 10709
rect 57513 10706 57579 10709
rect 56466 10704 57579 10706
rect 56466 10648 56598 10704
rect 56654 10648 57518 10704
rect 57574 10648 57579 10704
rect 56466 10646 57579 10648
rect 56550 10643 56659 10646
rect 57513 10643 57579 10646
rect 29269 10570 29335 10573
rect 30097 10570 30163 10573
rect 29269 10568 30163 10570
rect 29269 10512 29274 10568
rect 29330 10512 30102 10568
rect 30158 10512 30163 10568
rect 29269 10510 30163 10512
rect 29269 10507 29335 10510
rect 30097 10507 30163 10510
rect 30925 10570 30991 10573
rect 34237 10570 34303 10573
rect 30925 10568 34303 10570
rect 30925 10512 30930 10568
rect 30986 10512 34242 10568
rect 34298 10512 34303 10568
rect 30925 10510 34303 10512
rect 30925 10507 30991 10510
rect 34237 10507 34303 10510
rect 52177 10570 52243 10573
rect 56550 10570 56610 10643
rect 52177 10568 56610 10570
rect 52177 10512 52182 10568
rect 52238 10512 56610 10568
rect 52177 10510 56610 10512
rect 52177 10507 52243 10510
rect 26601 10434 26667 10437
rect 28533 10434 28599 10437
rect 26601 10432 28599 10434
rect 26601 10376 26606 10432
rect 26662 10376 28538 10432
rect 28594 10376 28599 10432
rect 26601 10374 28599 10376
rect 26601 10371 26667 10374
rect 28533 10371 28599 10374
rect 49509 10434 49575 10437
rect 49785 10434 49851 10437
rect 54661 10434 54727 10437
rect 49509 10432 54727 10434
rect 49509 10376 49514 10432
rect 49570 10376 49790 10432
rect 49846 10376 54666 10432
rect 54722 10376 54727 10432
rect 49509 10374 54727 10376
rect 49509 10371 49575 10374
rect 49785 10371 49851 10374
rect 54661 10371 54727 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 27470 10236 27476 10300
rect 27540 10298 27546 10300
rect 28441 10298 28507 10301
rect 34145 10298 34211 10301
rect 27540 10296 28507 10298
rect 27540 10240 28446 10296
rect 28502 10240 28507 10296
rect 27540 10238 28507 10240
rect 27540 10236 27546 10238
rect 28441 10235 28507 10238
rect 34102 10296 34211 10298
rect 34102 10240 34150 10296
rect 34206 10240 34211 10296
rect 34102 10235 34211 10240
rect 45921 10298 45987 10301
rect 46054 10298 46060 10300
rect 45921 10296 46060 10298
rect 45921 10240 45926 10296
rect 45982 10240 46060 10296
rect 45921 10238 46060 10240
rect 45921 10235 45987 10238
rect 46054 10236 46060 10238
rect 46124 10236 46130 10300
rect 27429 10162 27495 10165
rect 28257 10162 28323 10165
rect 29913 10162 29979 10165
rect 30925 10162 30991 10165
rect 31753 10162 31819 10165
rect 27429 10160 31819 10162
rect 27429 10104 27434 10160
rect 27490 10104 28262 10160
rect 28318 10104 29918 10160
rect 29974 10104 30930 10160
rect 30986 10104 31758 10160
rect 31814 10104 31819 10160
rect 27429 10102 31819 10104
rect 27429 10099 27495 10102
rect 28257 10099 28323 10102
rect 29913 10099 29979 10102
rect 30925 10099 30991 10102
rect 31753 10099 31819 10102
rect 31201 10026 31267 10029
rect 33685 10026 33751 10029
rect 31201 10024 33751 10026
rect 31201 9968 31206 10024
rect 31262 9968 33690 10024
rect 33746 9968 33751 10024
rect 31201 9966 33751 9968
rect 31201 9963 31267 9966
rect 33685 9963 33751 9966
rect 34102 9893 34162 10235
rect 46841 10162 46907 10165
rect 47342 10162 47348 10164
rect 46841 10160 47348 10162
rect 46841 10104 46846 10160
rect 46902 10104 47348 10160
rect 46841 10102 47348 10104
rect 46841 10099 46907 10102
rect 47342 10100 47348 10102
rect 47412 10162 47418 10164
rect 48773 10162 48839 10165
rect 47412 10160 48839 10162
rect 47412 10104 48778 10160
rect 48834 10104 48839 10160
rect 47412 10102 48839 10104
rect 47412 10100 47418 10102
rect 48773 10099 48839 10102
rect 41321 10026 41387 10029
rect 45277 10026 45343 10029
rect 41321 10024 45343 10026
rect 41321 9968 41326 10024
rect 41382 9968 45282 10024
rect 45338 9968 45343 10024
rect 41321 9966 45343 9968
rect 41321 9963 41387 9966
rect 45277 9963 45343 9966
rect 48589 10026 48655 10029
rect 49417 10026 49483 10029
rect 53649 10026 53715 10029
rect 48589 10024 53715 10026
rect 48589 9968 48594 10024
rect 48650 9968 49422 10024
rect 49478 9968 53654 10024
rect 53710 9968 53715 10024
rect 48589 9966 53715 9968
rect 48589 9963 48655 9966
rect 49417 9963 49483 9966
rect 53649 9963 53715 9966
rect 26325 9890 26391 9893
rect 28073 9890 28139 9893
rect 26325 9888 28139 9890
rect 26325 9832 26330 9888
rect 26386 9832 28078 9888
rect 28134 9832 28139 9888
rect 26325 9830 28139 9832
rect 34102 9888 34211 9893
rect 34102 9832 34150 9888
rect 34206 9832 34211 9888
rect 34102 9830 34211 9832
rect 26325 9827 26391 9830
rect 28073 9827 28139 9830
rect 34145 9827 34211 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 27613 9754 27679 9757
rect 32949 9754 33015 9757
rect 33317 9754 33383 9757
rect 27613 9752 33383 9754
rect 27613 9696 27618 9752
rect 27674 9696 32954 9752
rect 33010 9696 33322 9752
rect 33378 9696 33383 9752
rect 27613 9694 33383 9696
rect 27613 9691 27679 9694
rect 32949 9691 33015 9694
rect 33317 9691 33383 9694
rect 33910 9692 33916 9756
rect 33980 9754 33986 9756
rect 34053 9754 34119 9757
rect 33980 9752 34119 9754
rect 33980 9696 34058 9752
rect 34114 9696 34119 9752
rect 33980 9694 34119 9696
rect 33980 9692 33986 9694
rect 34053 9691 34119 9694
rect 43345 9754 43411 9757
rect 44357 9754 44423 9757
rect 43345 9752 44423 9754
rect 43345 9696 43350 9752
rect 43406 9696 44362 9752
rect 44418 9696 44423 9752
rect 43345 9694 44423 9696
rect 43345 9691 43411 9694
rect 44357 9691 44423 9694
rect 52453 9754 52519 9757
rect 53465 9754 53531 9757
rect 57237 9754 57303 9757
rect 52453 9752 57303 9754
rect 52453 9696 52458 9752
rect 52514 9696 53470 9752
rect 53526 9696 57242 9752
rect 57298 9696 57303 9752
rect 52453 9694 57303 9696
rect 52453 9691 52519 9694
rect 53465 9691 53531 9694
rect 57237 9691 57303 9694
rect 29177 9618 29243 9621
rect 29821 9620 29887 9621
rect 29821 9618 29868 9620
rect 29177 9616 29868 9618
rect 29177 9560 29182 9616
rect 29238 9560 29826 9616
rect 29177 9558 29868 9560
rect 29177 9555 29243 9558
rect 29821 9556 29868 9558
rect 29932 9556 29938 9620
rect 32121 9618 32187 9621
rect 41321 9618 41387 9621
rect 32121 9616 41387 9618
rect 32121 9560 32126 9616
rect 32182 9560 41326 9616
rect 41382 9560 41387 9616
rect 32121 9558 41387 9560
rect 29821 9555 29887 9556
rect 32121 9555 32187 9558
rect 41321 9555 41387 9558
rect 45829 9618 45895 9621
rect 52177 9618 52243 9621
rect 45829 9616 52243 9618
rect 45829 9560 45834 9616
rect 45890 9560 52182 9616
rect 52238 9560 52243 9616
rect 45829 9558 52243 9560
rect 45829 9555 45895 9558
rect 52177 9555 52243 9558
rect 52453 9618 52519 9621
rect 53741 9618 53807 9621
rect 52453 9616 53807 9618
rect 52453 9560 52458 9616
rect 52514 9560 53746 9616
rect 53802 9560 53807 9616
rect 52453 9558 53807 9560
rect 52453 9555 52519 9558
rect 53741 9555 53807 9558
rect 32305 9482 32371 9485
rect 33041 9482 33107 9485
rect 35801 9482 35867 9485
rect 32305 9480 35867 9482
rect 32305 9424 32310 9480
rect 32366 9424 33046 9480
rect 33102 9424 35806 9480
rect 35862 9424 35867 9480
rect 32305 9422 35867 9424
rect 32305 9419 32371 9422
rect 33041 9419 33107 9422
rect 35801 9419 35867 9422
rect 37273 9482 37339 9485
rect 38193 9482 38259 9485
rect 37273 9480 38259 9482
rect 37273 9424 37278 9480
rect 37334 9424 38198 9480
rect 38254 9424 38259 9480
rect 37273 9422 38259 9424
rect 37273 9419 37339 9422
rect 38193 9419 38259 9422
rect 43713 9482 43779 9485
rect 46289 9482 46355 9485
rect 43713 9480 46355 9482
rect 43713 9424 43718 9480
rect 43774 9424 46294 9480
rect 46350 9424 46355 9480
rect 43713 9422 46355 9424
rect 43713 9419 43779 9422
rect 46289 9419 46355 9422
rect 48497 9482 48563 9485
rect 51533 9482 51599 9485
rect 48497 9480 51599 9482
rect 48497 9424 48502 9480
rect 48558 9424 51538 9480
rect 51594 9424 51599 9480
rect 48497 9422 51599 9424
rect 48497 9419 48563 9422
rect 51533 9419 51599 9422
rect 36813 9346 36879 9349
rect 37641 9346 37707 9349
rect 36813 9344 37707 9346
rect 36813 9288 36818 9344
rect 36874 9288 37646 9344
rect 37702 9288 37707 9344
rect 36813 9286 37707 9288
rect 36813 9283 36879 9286
rect 37641 9283 37707 9286
rect 44817 9346 44883 9349
rect 47393 9346 47459 9349
rect 44817 9344 47459 9346
rect 44817 9288 44822 9344
rect 44878 9288 47398 9344
rect 47454 9288 47459 9344
rect 44817 9286 47459 9288
rect 44817 9283 44883 9286
rect 47393 9283 47459 9286
rect 48681 9346 48747 9349
rect 52545 9346 52611 9349
rect 48681 9344 52611 9346
rect 48681 9288 48686 9344
rect 48742 9288 52550 9344
rect 52606 9288 52611 9344
rect 48681 9286 52611 9288
rect 48681 9283 48747 9286
rect 52545 9283 52611 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 28901 9210 28967 9213
rect 30005 9210 30071 9213
rect 38837 9212 38903 9213
rect 38837 9210 38884 9212
rect 28901 9208 30071 9210
rect 28901 9152 28906 9208
rect 28962 9152 30010 9208
rect 30066 9152 30071 9208
rect 28901 9150 30071 9152
rect 38792 9208 38884 9210
rect 38792 9152 38842 9208
rect 38792 9150 38884 9152
rect 28901 9147 28967 9150
rect 30005 9147 30071 9150
rect 38837 9148 38884 9150
rect 38948 9148 38954 9212
rect 48957 9210 49023 9213
rect 50061 9210 50127 9213
rect 48957 9208 50127 9210
rect 48957 9152 48962 9208
rect 49018 9152 50066 9208
rect 50122 9152 50127 9208
rect 48957 9150 50127 9152
rect 38837 9147 38903 9148
rect 48957 9147 49023 9150
rect 50061 9147 50127 9150
rect 25405 9074 25471 9077
rect 28257 9074 28323 9077
rect 25405 9072 28323 9074
rect 25405 9016 25410 9072
rect 25466 9016 28262 9072
rect 28318 9016 28323 9072
rect 25405 9014 28323 9016
rect 25405 9011 25471 9014
rect 28257 9011 28323 9014
rect 29085 9074 29151 9077
rect 30005 9074 30071 9077
rect 29085 9072 30071 9074
rect 29085 9016 29090 9072
rect 29146 9016 30010 9072
rect 30066 9016 30071 9072
rect 29085 9014 30071 9016
rect 29085 9011 29151 9014
rect 30005 9011 30071 9014
rect 46289 9074 46355 9077
rect 47025 9074 47091 9077
rect 46289 9072 47091 9074
rect 46289 9016 46294 9072
rect 46350 9016 47030 9072
rect 47086 9016 47091 9072
rect 46289 9014 47091 9016
rect 46289 9011 46355 9014
rect 47025 9011 47091 9014
rect 27613 8938 27679 8941
rect 29637 8938 29703 8941
rect 27613 8936 29703 8938
rect 27613 8880 27618 8936
rect 27674 8880 29642 8936
rect 29698 8880 29703 8936
rect 27613 8878 29703 8880
rect 27613 8875 27679 8878
rect 29637 8875 29703 8878
rect 29821 8938 29887 8941
rect 32305 8938 32371 8941
rect 29821 8936 32371 8938
rect 29821 8880 29826 8936
rect 29882 8880 32310 8936
rect 32366 8880 32371 8936
rect 29821 8878 32371 8880
rect 29821 8875 29887 8878
rect 32305 8875 32371 8878
rect 32489 8938 32555 8941
rect 36169 8938 36235 8941
rect 32489 8936 36235 8938
rect 32489 8880 32494 8936
rect 32550 8880 36174 8936
rect 36230 8880 36235 8936
rect 32489 8878 36235 8880
rect 32489 8875 32555 8878
rect 36169 8875 36235 8878
rect 45645 8938 45711 8941
rect 46013 8938 46079 8941
rect 47301 8938 47367 8941
rect 47577 8938 47643 8941
rect 45645 8936 47643 8938
rect 45645 8880 45650 8936
rect 45706 8880 46018 8936
rect 46074 8880 47306 8936
rect 47362 8880 47582 8936
rect 47638 8880 47643 8936
rect 45645 8878 47643 8880
rect 45645 8875 45711 8878
rect 46013 8875 46079 8878
rect 47301 8875 47367 8878
rect 47577 8875 47643 8878
rect 51942 8876 51948 8940
rect 52012 8938 52018 8940
rect 52545 8938 52611 8941
rect 56409 8938 56475 8941
rect 52012 8936 56475 8938
rect 52012 8880 52550 8936
rect 52606 8880 56414 8936
rect 56470 8880 56475 8936
rect 52012 8878 56475 8880
rect 52012 8876 52018 8878
rect 52545 8875 52611 8878
rect 56409 8875 56475 8878
rect 27889 8802 27955 8805
rect 30925 8802 30991 8805
rect 27889 8800 30991 8802
rect 27889 8744 27894 8800
rect 27950 8744 30930 8800
rect 30986 8744 30991 8800
rect 27889 8742 30991 8744
rect 27889 8739 27955 8742
rect 30925 8739 30991 8742
rect 32765 8802 32831 8805
rect 35893 8802 35959 8805
rect 45645 8804 45711 8805
rect 45645 8802 45692 8804
rect 32765 8800 35959 8802
rect 32765 8744 32770 8800
rect 32826 8744 35898 8800
rect 35954 8744 35959 8800
rect 32765 8742 35959 8744
rect 45600 8800 45692 8802
rect 45600 8744 45650 8800
rect 45600 8742 45692 8744
rect 32765 8739 32831 8742
rect 35893 8739 35959 8742
rect 45645 8740 45692 8742
rect 45756 8740 45762 8804
rect 45645 8739 45711 8740
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 30281 8666 30347 8669
rect 30281 8664 33978 8666
rect 30281 8608 30286 8664
rect 30342 8608 33978 8664
rect 30281 8606 33978 8608
rect 30281 8603 30347 8606
rect 31385 8530 31451 8533
rect 32121 8530 32187 8533
rect 31385 8528 32187 8530
rect 31385 8472 31390 8528
rect 31446 8472 32126 8528
rect 32182 8472 32187 8528
rect 31385 8470 32187 8472
rect 33918 8530 33978 8606
rect 35249 8530 35315 8533
rect 33918 8528 35315 8530
rect 33918 8472 35254 8528
rect 35310 8472 35315 8528
rect 33918 8470 35315 8472
rect 31385 8467 31451 8470
rect 32121 8467 32187 8470
rect 35249 8467 35315 8470
rect 45369 8530 45435 8533
rect 48313 8530 48379 8533
rect 45369 8528 48379 8530
rect 45369 8472 45374 8528
rect 45430 8472 48318 8528
rect 48374 8472 48379 8528
rect 45369 8470 48379 8472
rect 45369 8467 45435 8470
rect 48313 8467 48379 8470
rect 49601 8530 49667 8533
rect 50613 8530 50679 8533
rect 51349 8530 51415 8533
rect 49601 8528 51415 8530
rect 49601 8472 49606 8528
rect 49662 8472 50618 8528
rect 50674 8472 51354 8528
rect 51410 8472 51415 8528
rect 49601 8470 51415 8472
rect 49601 8467 49667 8470
rect 50613 8467 50679 8470
rect 51349 8467 51415 8470
rect 29310 8332 29316 8396
rect 29380 8394 29386 8396
rect 29453 8394 29519 8397
rect 29380 8392 29519 8394
rect 29380 8336 29458 8392
rect 29514 8336 29519 8392
rect 29380 8334 29519 8336
rect 29380 8332 29386 8334
rect 29453 8331 29519 8334
rect 30281 8394 30347 8397
rect 37273 8394 37339 8397
rect 30281 8392 37339 8394
rect 30281 8336 30286 8392
rect 30342 8336 37278 8392
rect 37334 8336 37339 8392
rect 30281 8334 37339 8336
rect 30281 8331 30347 8334
rect 37273 8331 37339 8334
rect 28022 8196 28028 8260
rect 28092 8258 28098 8260
rect 32029 8258 32095 8261
rect 28092 8256 32095 8258
rect 28092 8200 32034 8256
rect 32090 8200 32095 8256
rect 28092 8198 32095 8200
rect 28092 8196 28098 8198
rect 32029 8195 32095 8198
rect 48313 8258 48379 8261
rect 49366 8258 49372 8260
rect 48313 8256 49372 8258
rect 48313 8200 48318 8256
rect 48374 8200 49372 8256
rect 48313 8198 49372 8200
rect 48313 8195 48379 8198
rect 49366 8196 49372 8198
rect 49436 8258 49442 8260
rect 54201 8258 54267 8261
rect 49436 8256 54267 8258
rect 49436 8200 54206 8256
rect 54262 8200 54267 8256
rect 49436 8198 54267 8200
rect 49436 8196 49442 8198
rect 54201 8195 54267 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 32765 8122 32831 8125
rect 34513 8122 34579 8125
rect 32765 8120 34579 8122
rect 32765 8064 32770 8120
rect 32826 8064 34518 8120
rect 34574 8064 34579 8120
rect 32765 8062 34579 8064
rect 32765 8059 32831 8062
rect 34513 8059 34579 8062
rect 51206 8060 51212 8124
rect 51276 8122 51282 8124
rect 51809 8122 51875 8125
rect 51276 8120 51875 8122
rect 51276 8064 51814 8120
rect 51870 8064 51875 8120
rect 51276 8062 51875 8064
rect 51276 8060 51282 8062
rect 51809 8059 51875 8062
rect 29085 7986 29151 7989
rect 30005 7986 30071 7989
rect 31753 7986 31819 7989
rect 29085 7984 31819 7986
rect 29085 7928 29090 7984
rect 29146 7928 30010 7984
rect 30066 7928 31758 7984
rect 31814 7928 31819 7984
rect 29085 7926 31819 7928
rect 29085 7923 29151 7926
rect 30005 7923 30071 7926
rect 31753 7923 31819 7926
rect 35157 7986 35223 7989
rect 35985 7986 36051 7989
rect 35157 7984 36051 7986
rect 35157 7928 35162 7984
rect 35218 7928 35990 7984
rect 36046 7928 36051 7984
rect 35157 7926 36051 7928
rect 35157 7923 35223 7926
rect 35985 7923 36051 7926
rect 34145 7850 34211 7853
rect 38377 7850 38443 7853
rect 34145 7848 38443 7850
rect 34145 7792 34150 7848
rect 34206 7792 38382 7848
rect 38438 7792 38443 7848
rect 34145 7790 38443 7792
rect 34145 7787 34211 7790
rect 38377 7787 38443 7790
rect 44541 7850 44607 7853
rect 47669 7850 47735 7853
rect 44541 7848 47735 7850
rect 44541 7792 44546 7848
rect 44602 7792 47674 7848
rect 47730 7792 47735 7848
rect 44541 7790 47735 7792
rect 44541 7787 44607 7790
rect 47669 7787 47735 7790
rect 29310 7652 29316 7716
rect 29380 7714 29386 7716
rect 29453 7714 29519 7717
rect 29380 7712 29519 7714
rect 29380 7656 29458 7712
rect 29514 7656 29519 7712
rect 29380 7654 29519 7656
rect 29380 7652 29386 7654
rect 29453 7651 29519 7654
rect 49325 7714 49391 7717
rect 49877 7714 49943 7717
rect 49325 7712 49943 7714
rect 49325 7656 49330 7712
rect 49386 7656 49882 7712
rect 49938 7656 49943 7712
rect 49325 7654 49943 7656
rect 49325 7651 49391 7654
rect 49877 7651 49943 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 31201 7578 31267 7581
rect 35617 7578 35683 7581
rect 31201 7576 35683 7578
rect 31201 7520 31206 7576
rect 31262 7520 35622 7576
rect 35678 7520 35683 7576
rect 31201 7518 35683 7520
rect 31201 7515 31267 7518
rect 35617 7515 35683 7518
rect 27613 7442 27679 7445
rect 27981 7442 28047 7445
rect 27613 7440 28047 7442
rect 27613 7384 27618 7440
rect 27674 7384 27986 7440
rect 28042 7384 28047 7440
rect 27613 7382 28047 7384
rect 27613 7379 27679 7382
rect 27981 7379 28047 7382
rect 30097 7442 30163 7445
rect 31109 7442 31175 7445
rect 30097 7440 31175 7442
rect 30097 7384 30102 7440
rect 30158 7384 31114 7440
rect 31170 7384 31175 7440
rect 30097 7382 31175 7384
rect 30097 7379 30163 7382
rect 31109 7379 31175 7382
rect 31661 7442 31727 7445
rect 32489 7442 32555 7445
rect 35934 7442 35940 7444
rect 31661 7440 35940 7442
rect 31661 7384 31666 7440
rect 31722 7384 32494 7440
rect 32550 7384 35940 7440
rect 31661 7382 35940 7384
rect 31661 7379 31727 7382
rect 32489 7379 32555 7382
rect 35934 7380 35940 7382
rect 36004 7380 36010 7444
rect 49601 7442 49667 7445
rect 55213 7442 55279 7445
rect 49601 7440 55279 7442
rect 49601 7384 49606 7440
rect 49662 7384 55218 7440
rect 55274 7384 55279 7440
rect 49601 7382 55279 7384
rect 49601 7379 49667 7382
rect 55213 7379 55279 7382
rect 26734 7244 26740 7308
rect 26804 7306 26810 7308
rect 27981 7306 28047 7309
rect 35525 7306 35591 7309
rect 26804 7304 28047 7306
rect 26804 7248 27986 7304
rect 28042 7248 28047 7304
rect 26804 7246 28047 7248
rect 26804 7244 26810 7246
rect 27981 7243 28047 7246
rect 34792 7304 35591 7306
rect 34792 7248 35530 7304
rect 35586 7248 35591 7304
rect 34792 7246 35591 7248
rect 33225 7170 33291 7173
rect 34792 7170 34852 7246
rect 35525 7243 35591 7246
rect 46749 7306 46815 7309
rect 51073 7306 51139 7309
rect 46749 7304 51139 7306
rect 46749 7248 46754 7304
rect 46810 7248 51078 7304
rect 51134 7248 51139 7304
rect 46749 7246 51139 7248
rect 46749 7243 46815 7246
rect 51073 7243 51139 7246
rect 43713 7172 43779 7173
rect 43662 7170 43668 7172
rect 33225 7168 34852 7170
rect 33225 7112 33230 7168
rect 33286 7112 34852 7168
rect 33225 7110 34852 7112
rect 43622 7110 43668 7170
rect 43732 7168 43779 7172
rect 43774 7112 43779 7168
rect 33225 7107 33291 7110
rect 43662 7108 43668 7110
rect 43732 7108 43779 7112
rect 43713 7107 43779 7108
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 27061 7034 27127 7037
rect 28349 7034 28415 7037
rect 27061 7032 28415 7034
rect 27061 6976 27066 7032
rect 27122 6976 28354 7032
rect 28410 6976 28415 7032
rect 27061 6974 28415 6976
rect 27061 6971 27127 6974
rect 28349 6971 28415 6974
rect 31661 7034 31727 7037
rect 31845 7034 31911 7037
rect 31661 7032 31911 7034
rect 31661 6976 31666 7032
rect 31722 6976 31850 7032
rect 31906 6976 31911 7032
rect 31661 6974 31911 6976
rect 31661 6971 31727 6974
rect 31845 6971 31911 6974
rect 48865 7034 48931 7037
rect 53373 7034 53439 7037
rect 48865 7032 53439 7034
rect 48865 6976 48870 7032
rect 48926 6976 53378 7032
rect 53434 6976 53439 7032
rect 48865 6974 53439 6976
rect 48865 6971 48931 6974
rect 53373 6971 53439 6974
rect 26785 6898 26851 6901
rect 29177 6898 29243 6901
rect 36077 6898 36143 6901
rect 36445 6898 36511 6901
rect 26785 6896 36511 6898
rect 26785 6840 26790 6896
rect 26846 6840 29182 6896
rect 29238 6840 36082 6896
rect 36138 6840 36450 6896
rect 36506 6840 36511 6896
rect 26785 6838 36511 6840
rect 26785 6835 26851 6838
rect 29177 6835 29243 6838
rect 36077 6835 36143 6838
rect 36445 6835 36511 6838
rect 43897 6898 43963 6901
rect 44582 6898 44588 6900
rect 43897 6896 44588 6898
rect 43897 6840 43902 6896
rect 43958 6840 44588 6896
rect 43897 6838 44588 6840
rect 43897 6835 43963 6838
rect 44582 6836 44588 6838
rect 44652 6836 44658 6900
rect 48313 6898 48379 6901
rect 48446 6898 48452 6900
rect 48313 6896 48452 6898
rect 48313 6840 48318 6896
rect 48374 6840 48452 6896
rect 48313 6838 48452 6840
rect 48313 6835 48379 6838
rect 48446 6836 48452 6838
rect 48516 6836 48522 6900
rect 57881 6898 57947 6901
rect 59200 6898 59800 6928
rect 57881 6896 59800 6898
rect 57881 6840 57886 6896
rect 57942 6840 59800 6896
rect 57881 6838 59800 6840
rect 57881 6835 57947 6838
rect 59200 6808 59800 6838
rect 31150 6700 31156 6764
rect 31220 6762 31226 6764
rect 32489 6762 32555 6765
rect 31220 6760 32555 6762
rect 31220 6704 32494 6760
rect 32550 6704 32555 6760
rect 31220 6702 32555 6704
rect 31220 6700 31226 6702
rect 32489 6699 32555 6702
rect 49785 6762 49851 6765
rect 50337 6762 50403 6765
rect 49785 6760 50403 6762
rect 49785 6704 49790 6760
rect 49846 6704 50342 6760
rect 50398 6704 50403 6760
rect 49785 6702 50403 6704
rect 49785 6699 49851 6702
rect 50337 6699 50403 6702
rect 54845 6762 54911 6765
rect 55070 6762 55076 6764
rect 54845 6760 55076 6762
rect 54845 6704 54850 6760
rect 54906 6704 55076 6760
rect 54845 6702 55076 6704
rect 54845 6699 54911 6702
rect 55070 6700 55076 6702
rect 55140 6700 55146 6764
rect 33501 6626 33567 6629
rect 33777 6626 33843 6629
rect 33501 6624 33843 6626
rect 33501 6568 33506 6624
rect 33562 6568 33782 6624
rect 33838 6568 33843 6624
rect 33501 6566 33843 6568
rect 33501 6563 33567 6566
rect 33777 6563 33843 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 29821 6490 29887 6493
rect 32121 6490 32187 6493
rect 37917 6490 37983 6493
rect 29821 6488 37983 6490
rect 29821 6432 29826 6488
rect 29882 6432 32126 6488
rect 32182 6432 37922 6488
rect 37978 6432 37983 6488
rect 29821 6430 37983 6432
rect 29821 6427 29887 6430
rect 32121 6427 32187 6430
rect 37917 6427 37983 6430
rect 38653 6354 38719 6357
rect 40401 6354 40467 6357
rect 38653 6352 40467 6354
rect 38653 6296 38658 6352
rect 38714 6296 40406 6352
rect 40462 6296 40467 6352
rect 38653 6294 40467 6296
rect 38653 6291 38719 6294
rect 40401 6291 40467 6294
rect 47669 6354 47735 6357
rect 50337 6354 50403 6357
rect 47669 6352 50403 6354
rect 47669 6296 47674 6352
rect 47730 6296 50342 6352
rect 50398 6296 50403 6352
rect 47669 6294 50403 6296
rect 47669 6291 47735 6294
rect 50337 6291 50403 6294
rect 51165 6354 51231 6357
rect 51717 6354 51783 6357
rect 51165 6352 51783 6354
rect 51165 6296 51170 6352
rect 51226 6296 51722 6352
rect 51778 6296 51783 6352
rect 51165 6294 51783 6296
rect 51165 6291 51231 6294
rect 51717 6291 51783 6294
rect 27337 6218 27403 6221
rect 32581 6218 32647 6221
rect 34145 6218 34211 6221
rect 27337 6216 34211 6218
rect 27337 6160 27342 6216
rect 27398 6160 32586 6216
rect 32642 6160 34150 6216
rect 34206 6160 34211 6216
rect 27337 6158 34211 6160
rect 27337 6155 27403 6158
rect 32581 6155 32647 6158
rect 34145 6155 34211 6158
rect 28717 6082 28783 6085
rect 29269 6082 29335 6085
rect 31385 6082 31451 6085
rect 28717 6080 31451 6082
rect 28717 6024 28722 6080
rect 28778 6024 29274 6080
rect 29330 6024 31390 6080
rect 31446 6024 31451 6080
rect 28717 6022 31451 6024
rect 28717 6019 28783 6022
rect 29269 6019 29335 6022
rect 31385 6019 31451 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 31385 5946 31451 5949
rect 31518 5946 31524 5948
rect 31385 5944 31524 5946
rect 31385 5888 31390 5944
rect 31446 5888 31524 5944
rect 31385 5886 31524 5888
rect 31385 5883 31451 5886
rect 31518 5884 31524 5886
rect 31588 5884 31594 5948
rect 38285 5810 38351 5813
rect 39798 5810 39804 5812
rect 38285 5808 39804 5810
rect 38285 5752 38290 5808
rect 38346 5752 39804 5808
rect 38285 5750 39804 5752
rect 38285 5747 38351 5750
rect 39798 5748 39804 5750
rect 39868 5748 39874 5812
rect 43253 5810 43319 5813
rect 49601 5810 49667 5813
rect 43253 5808 49667 5810
rect 43253 5752 43258 5808
rect 43314 5752 49606 5808
rect 49662 5752 49667 5808
rect 43253 5750 49667 5752
rect 43253 5747 43319 5750
rect 49601 5747 49667 5750
rect 22645 5674 22711 5677
rect 29913 5674 29979 5677
rect 22645 5672 29979 5674
rect 22645 5616 22650 5672
rect 22706 5616 29918 5672
rect 29974 5616 29979 5672
rect 22645 5614 29979 5616
rect 22645 5611 22711 5614
rect 29913 5611 29979 5614
rect 46013 5674 46079 5677
rect 49693 5674 49759 5677
rect 46013 5672 49759 5674
rect 46013 5616 46018 5672
rect 46074 5616 49698 5672
rect 49754 5616 49759 5672
rect 46013 5614 49759 5616
rect 46013 5611 46079 5614
rect 49693 5611 49759 5614
rect 200 5538 800 5568
rect 1669 5538 1735 5541
rect 200 5536 1735 5538
rect 200 5480 1674 5536
rect 1730 5480 1735 5536
rect 200 5478 1735 5480
rect 200 5448 800 5478
rect 1669 5475 1735 5478
rect 26049 5538 26115 5541
rect 28441 5538 28507 5541
rect 28901 5538 28967 5541
rect 26049 5536 28967 5538
rect 26049 5480 26054 5536
rect 26110 5480 28446 5536
rect 28502 5480 28906 5536
rect 28962 5480 28967 5536
rect 26049 5478 28967 5480
rect 26049 5475 26115 5478
rect 28441 5475 28507 5478
rect 28901 5475 28967 5478
rect 37273 5538 37339 5541
rect 37590 5538 37596 5540
rect 37273 5536 37596 5538
rect 37273 5480 37278 5536
rect 37334 5480 37596 5536
rect 37273 5478 37596 5480
rect 37273 5475 37339 5478
rect 37590 5476 37596 5478
rect 37660 5538 37666 5540
rect 37825 5538 37891 5541
rect 37660 5536 37891 5538
rect 37660 5480 37830 5536
rect 37886 5480 37891 5536
rect 37660 5478 37891 5480
rect 37660 5476 37666 5478
rect 37825 5475 37891 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 27613 5402 27679 5405
rect 28717 5402 28783 5405
rect 27613 5400 28783 5402
rect 27613 5344 27618 5400
rect 27674 5344 28722 5400
rect 28778 5344 28783 5400
rect 27613 5342 28783 5344
rect 27613 5339 27679 5342
rect 28717 5339 28783 5342
rect 30097 5402 30163 5405
rect 30230 5402 30236 5404
rect 30097 5400 30236 5402
rect 30097 5344 30102 5400
rect 30158 5344 30236 5400
rect 30097 5342 30236 5344
rect 30097 5339 30163 5342
rect 30230 5340 30236 5342
rect 30300 5340 30306 5404
rect 33777 5402 33843 5405
rect 33910 5402 33916 5404
rect 33777 5400 33916 5402
rect 33777 5344 33782 5400
rect 33838 5344 33916 5400
rect 33777 5342 33916 5344
rect 33777 5339 33843 5342
rect 33910 5340 33916 5342
rect 33980 5340 33986 5404
rect 35065 5402 35131 5405
rect 38009 5402 38075 5405
rect 35065 5400 38075 5402
rect 35065 5344 35070 5400
rect 35126 5344 38014 5400
rect 38070 5344 38075 5400
rect 35065 5342 38075 5344
rect 35065 5339 35131 5342
rect 38009 5339 38075 5342
rect 1761 5266 1827 5269
rect 41413 5266 41479 5269
rect 1761 5264 41479 5266
rect 1761 5208 1766 5264
rect 1822 5208 41418 5264
rect 41474 5208 41479 5264
rect 1761 5206 41479 5208
rect 1761 5203 1827 5206
rect 41413 5203 41479 5206
rect 46565 5266 46631 5269
rect 51533 5266 51599 5269
rect 51942 5266 51948 5268
rect 46565 5264 51948 5266
rect 46565 5208 46570 5264
rect 46626 5208 51538 5264
rect 51594 5208 51948 5264
rect 46565 5206 51948 5208
rect 46565 5203 46631 5206
rect 51533 5203 51599 5206
rect 51942 5204 51948 5206
rect 52012 5204 52018 5268
rect 28533 5130 28599 5133
rect 34329 5130 34395 5133
rect 35709 5130 35775 5133
rect 28533 5128 35775 5130
rect 28533 5072 28538 5128
rect 28594 5072 34334 5128
rect 34390 5072 35714 5128
rect 35770 5072 35775 5128
rect 28533 5070 35775 5072
rect 28533 5067 28599 5070
rect 34329 5067 34395 5070
rect 35709 5067 35775 5070
rect 46381 5130 46447 5133
rect 48497 5130 48563 5133
rect 46381 5128 48563 5130
rect 46381 5072 46386 5128
rect 46442 5072 48502 5128
rect 48558 5072 48563 5128
rect 46381 5070 48563 5072
rect 46381 5067 46447 5070
rect 48497 5067 48563 5070
rect 28625 4994 28691 4997
rect 33869 4994 33935 4997
rect 28625 4992 33935 4994
rect 28625 4936 28630 4992
rect 28686 4936 33874 4992
rect 33930 4936 33935 4992
rect 28625 4934 33935 4936
rect 28625 4931 28691 4934
rect 33869 4931 33935 4934
rect 47025 4994 47091 4997
rect 47669 4994 47735 4997
rect 47025 4992 47735 4994
rect 47025 4936 47030 4992
rect 47086 4936 47674 4992
rect 47730 4936 47735 4992
rect 47025 4934 47735 4936
rect 47025 4931 47091 4934
rect 47669 4931 47735 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 45185 4858 45251 4861
rect 47393 4858 47459 4861
rect 45185 4856 47459 4858
rect 45185 4800 45190 4856
rect 45246 4800 47398 4856
rect 47454 4800 47459 4856
rect 45185 4798 47459 4800
rect 45185 4795 45251 4798
rect 47393 4795 47459 4798
rect 42149 4722 42215 4725
rect 44449 4722 44515 4725
rect 46657 4722 46723 4725
rect 42149 4720 46723 4722
rect 42149 4664 42154 4720
rect 42210 4664 44454 4720
rect 44510 4664 46662 4720
rect 46718 4664 46723 4720
rect 42149 4662 46723 4664
rect 42149 4659 42215 4662
rect 44449 4659 44515 4662
rect 46657 4659 46723 4662
rect 36077 4586 36143 4589
rect 51625 4586 51691 4589
rect 36077 4584 51691 4586
rect 36077 4528 36082 4584
rect 36138 4528 51630 4584
rect 51686 4528 51691 4584
rect 36077 4526 51691 4528
rect 36077 4523 36143 4526
rect 51625 4523 51691 4526
rect 47577 4450 47643 4453
rect 47945 4450 48011 4453
rect 47577 4448 48011 4450
rect 47577 4392 47582 4448
rect 47638 4392 47950 4448
rect 48006 4392 48011 4448
rect 47577 4390 48011 4392
rect 47577 4387 47643 4390
rect 47945 4387 48011 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 27838 3980 27844 4044
rect 27908 4042 27914 4044
rect 27981 4042 28047 4045
rect 27908 4040 28047 4042
rect 27908 3984 27986 4040
rect 28042 3984 28047 4040
rect 27908 3982 28047 3984
rect 27908 3980 27914 3982
rect 27981 3979 28047 3982
rect 36118 3980 36124 4044
rect 36188 4042 36194 4044
rect 41505 4042 41571 4045
rect 36188 4040 41571 4042
rect 36188 3984 41510 4040
rect 41566 3984 41571 4040
rect 36188 3982 41571 3984
rect 36188 3980 36194 3982
rect 41505 3979 41571 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 47025 2682 47091 2685
rect 49918 2682 49924 2684
rect 47025 2680 49924 2682
rect 47025 2624 47030 2680
rect 47086 2624 49924 2680
rect 47025 2622 49924 2624
rect 47025 2619 47091 2622
rect 49918 2620 49924 2622
rect 49988 2620 49994 2684
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 59200 778 59800 808
rect 59905 778 59971 781
rect 59200 776 59971 778
rect 59200 720 59910 776
rect 59966 720 59971 776
rect 59200 718 59971 720
rect 59200 688 59800 718
rect 59905 715 59971 718
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 28028 57216 28092 57220
rect 28028 57160 28042 57216
rect 28042 57160 28092 57216
rect 28028 57156 28092 57160
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 49924 27644 49988 27708
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 49372 24788 49436 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 46060 22536 46124 22540
rect 46060 22480 46110 22536
rect 46110 22480 46124 22536
rect 46060 22476 46124 22480
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 53420 21252 53484 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 49188 20904 49252 20908
rect 49188 20848 49202 20904
rect 49202 20848 49252 20904
rect 49188 20844 49252 20848
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 44588 20300 44652 20364
rect 36124 20224 36188 20228
rect 36124 20168 36138 20224
rect 36138 20168 36188 20224
rect 36124 20164 36188 20168
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 43668 19408 43732 19412
rect 43668 19352 43682 19408
rect 43682 19352 43732 19408
rect 43668 19348 43732 19352
rect 52316 19212 52380 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 44036 17988 44100 18052
rect 53972 18048 54036 18052
rect 53972 17992 54022 18048
rect 54022 17992 54036 18048
rect 53972 17988 54036 17992
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 45692 17776 45756 17780
rect 45692 17720 45742 17776
rect 45742 17720 45756 17776
rect 45692 17716 45756 17720
rect 27476 17640 27540 17644
rect 27476 17584 27526 17640
rect 27526 17584 27540 17640
rect 27476 17580 27540 17584
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 38884 17096 38948 17100
rect 38884 17040 38934 17096
rect 38934 17040 38948 17096
rect 38884 17036 38948 17040
rect 48268 17096 48332 17100
rect 48268 17040 48318 17096
rect 48318 17040 48332 17096
rect 48268 17036 48332 17040
rect 48636 17036 48700 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 31524 16688 31588 16692
rect 31524 16632 31574 16688
rect 31574 16632 31588 16688
rect 31524 16628 31588 16632
rect 53788 16628 53852 16692
rect 49188 16492 49252 16556
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 45324 15464 45388 15468
rect 45324 15408 45374 15464
rect 45374 15408 45388 15464
rect 45324 15404 45388 15408
rect 49188 15464 49252 15468
rect 49188 15408 49238 15464
rect 49238 15408 49252 15464
rect 49188 15404 49252 15408
rect 30236 15268 30300 15332
rect 45508 15268 45572 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 53420 15132 53484 15196
rect 49372 14920 49436 14924
rect 49372 14864 49386 14920
rect 49386 14864 49436 14920
rect 49372 14860 49436 14864
rect 48636 14724 48700 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 31156 13772 31220 13836
rect 39804 13832 39868 13836
rect 39804 13776 39854 13832
rect 39854 13776 39868 13832
rect 39804 13772 39868 13776
rect 49372 13636 49436 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 48452 13560 48516 13564
rect 48452 13504 48502 13560
rect 48502 13504 48516 13560
rect 48452 13500 48516 13504
rect 48636 13288 48700 13292
rect 48636 13232 48650 13288
rect 48650 13232 48700 13288
rect 48636 13228 48700 13232
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 47348 13092 47412 13156
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 45508 12820 45572 12884
rect 50844 12820 50908 12884
rect 49188 12548 49252 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 52316 12276 52380 12340
rect 53788 12276 53852 12340
rect 29868 12140 29932 12204
rect 37596 12200 37660 12204
rect 37596 12144 37646 12200
rect 37646 12144 37660 12200
rect 37596 12140 37660 12144
rect 48268 12140 48332 12204
rect 26740 12004 26804 12068
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 44036 11868 44100 11932
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 27844 11052 27908 11116
rect 35940 11052 36004 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 45324 10780 45388 10844
rect 53972 10840 54036 10844
rect 53972 10784 54022 10840
rect 54022 10784 54036 10840
rect 53972 10780 54036 10784
rect 55076 10840 55140 10844
rect 55076 10784 55126 10840
rect 55126 10784 55140 10840
rect 55076 10780 55140 10784
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 27476 10236 27540 10300
rect 46060 10236 46124 10300
rect 47348 10100 47412 10164
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 33916 9692 33980 9756
rect 29868 9616 29932 9620
rect 29868 9560 29882 9616
rect 29882 9560 29932 9616
rect 29868 9556 29932 9560
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 38884 9208 38948 9212
rect 38884 9152 38898 9208
rect 38898 9152 38948 9208
rect 38884 9148 38948 9152
rect 51948 8876 52012 8940
rect 45692 8800 45756 8804
rect 45692 8744 45706 8800
rect 45706 8744 45756 8800
rect 45692 8740 45756 8744
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 29316 8332 29380 8396
rect 28028 8196 28092 8260
rect 49372 8196 49436 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 51212 8060 51276 8124
rect 29316 7652 29380 7716
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 35940 7380 36004 7444
rect 26740 7244 26804 7308
rect 43668 7168 43732 7172
rect 43668 7112 43718 7168
rect 43718 7112 43732 7168
rect 43668 7108 43732 7112
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 44588 6836 44652 6900
rect 48452 6836 48516 6900
rect 31156 6700 31220 6764
rect 55076 6700 55140 6764
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 31524 5884 31588 5948
rect 39804 5748 39868 5812
rect 37596 5476 37660 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 30236 5340 30300 5404
rect 33916 5340 33980 5404
rect 51948 5204 52012 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 27844 3980 27908 4044
rect 36124 3980 36188 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 49924 2620 49988 2684
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 28027 57220 28093 57221
rect 28027 57156 28028 57220
rect 28092 57156 28093 57220
rect 28027 57155 28093 57156
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 27475 17644 27541 17645
rect 27475 17580 27476 17644
rect 27540 17580 27541 17644
rect 27475 17579 27541 17580
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 26739 12068 26805 12069
rect 26739 12004 26740 12068
rect 26804 12004 26805 12068
rect 26739 12003 26805 12004
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 26742 7309 26802 12003
rect 27478 10301 27538 17579
rect 27843 11116 27909 11117
rect 27843 11052 27844 11116
rect 27908 11052 27909 11116
rect 27843 11051 27909 11052
rect 27475 10300 27541 10301
rect 27475 10236 27476 10300
rect 27540 10236 27541 10300
rect 27475 10235 27541 10236
rect 26739 7308 26805 7309
rect 26739 7244 26740 7308
rect 26804 7244 26805 7308
rect 26739 7243 26805 7244
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 27846 4045 27906 11051
rect 28030 8261 28090 57155
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 49923 27708 49989 27709
rect 49923 27644 49924 27708
rect 49988 27644 49989 27708
rect 49923 27643 49989 27644
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 49371 24852 49437 24853
rect 49371 24788 49372 24852
rect 49436 24788 49437 24852
rect 49371 24787 49437 24788
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 46059 22540 46125 22541
rect 46059 22476 46060 22540
rect 46124 22476 46125 22540
rect 46059 22475 46125 22476
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 44587 20364 44653 20365
rect 44587 20300 44588 20364
rect 44652 20300 44653 20364
rect 44587 20299 44653 20300
rect 36123 20228 36189 20229
rect 36123 20164 36124 20228
rect 36188 20164 36189 20228
rect 36123 20163 36189 20164
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 31523 16692 31589 16693
rect 31523 16628 31524 16692
rect 31588 16628 31589 16692
rect 31523 16627 31589 16628
rect 30235 15332 30301 15333
rect 30235 15268 30236 15332
rect 30300 15268 30301 15332
rect 30235 15267 30301 15268
rect 29867 12204 29933 12205
rect 29867 12140 29868 12204
rect 29932 12140 29933 12204
rect 29867 12139 29933 12140
rect 29870 9621 29930 12139
rect 29867 9620 29933 9621
rect 29867 9556 29868 9620
rect 29932 9556 29933 9620
rect 29867 9555 29933 9556
rect 29315 8396 29381 8397
rect 29315 8332 29316 8396
rect 29380 8332 29381 8396
rect 29315 8331 29381 8332
rect 28027 8260 28093 8261
rect 28027 8196 28028 8260
rect 28092 8196 28093 8260
rect 28027 8195 28093 8196
rect 29318 7717 29378 8331
rect 29315 7716 29381 7717
rect 29315 7652 29316 7716
rect 29380 7652 29381 7716
rect 29315 7651 29381 7652
rect 30238 5405 30298 15267
rect 31155 13836 31221 13837
rect 31155 13772 31156 13836
rect 31220 13772 31221 13836
rect 31155 13771 31221 13772
rect 31158 6765 31218 13771
rect 31155 6764 31221 6765
rect 31155 6700 31156 6764
rect 31220 6700 31221 6764
rect 31155 6699 31221 6700
rect 31526 5949 31586 16627
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 35939 11116 36005 11117
rect 35939 11052 35940 11116
rect 36004 11052 36005 11116
rect 35939 11051 36005 11052
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 33915 9756 33981 9757
rect 33915 9692 33916 9756
rect 33980 9692 33981 9756
rect 33915 9691 33981 9692
rect 31523 5948 31589 5949
rect 31523 5884 31524 5948
rect 31588 5884 31589 5948
rect 31523 5883 31589 5884
rect 33918 5405 33978 9691
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 35942 7445 36002 11051
rect 35939 7444 36005 7445
rect 35939 7380 35940 7444
rect 36004 7380 36005 7444
rect 35939 7379 36005 7380
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 30235 5404 30301 5405
rect 30235 5340 30236 5404
rect 30300 5340 30301 5404
rect 30235 5339 30301 5340
rect 33915 5404 33981 5405
rect 33915 5340 33916 5404
rect 33980 5340 33981 5404
rect 33915 5339 33981 5340
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 27843 4044 27909 4045
rect 27843 3980 27844 4044
rect 27908 3980 27909 4044
rect 27843 3979 27909 3980
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 3840 35248 4864
rect 36126 4045 36186 20163
rect 43667 19412 43733 19413
rect 43667 19348 43668 19412
rect 43732 19348 43733 19412
rect 43667 19347 43733 19348
rect 38883 17100 38949 17101
rect 38883 17036 38884 17100
rect 38948 17036 38949 17100
rect 38883 17035 38949 17036
rect 37595 12204 37661 12205
rect 37595 12140 37596 12204
rect 37660 12140 37661 12204
rect 37595 12139 37661 12140
rect 37598 5541 37658 12139
rect 38886 9213 38946 17035
rect 39803 13836 39869 13837
rect 39803 13772 39804 13836
rect 39868 13772 39869 13836
rect 39803 13771 39869 13772
rect 38883 9212 38949 9213
rect 38883 9148 38884 9212
rect 38948 9148 38949 9212
rect 38883 9147 38949 9148
rect 39806 5813 39866 13771
rect 43670 7173 43730 19347
rect 44035 18052 44101 18053
rect 44035 17988 44036 18052
rect 44100 17988 44101 18052
rect 44035 17987 44101 17988
rect 44038 11933 44098 17987
rect 44035 11932 44101 11933
rect 44035 11868 44036 11932
rect 44100 11868 44101 11932
rect 44035 11867 44101 11868
rect 43667 7172 43733 7173
rect 43667 7108 43668 7172
rect 43732 7108 43733 7172
rect 43667 7107 43733 7108
rect 44590 6901 44650 20299
rect 45691 17780 45757 17781
rect 45691 17716 45692 17780
rect 45756 17716 45757 17780
rect 45691 17715 45757 17716
rect 45323 15468 45389 15469
rect 45323 15404 45324 15468
rect 45388 15404 45389 15468
rect 45323 15403 45389 15404
rect 45326 10845 45386 15403
rect 45507 15332 45573 15333
rect 45507 15268 45508 15332
rect 45572 15268 45573 15332
rect 45507 15267 45573 15268
rect 45510 12885 45570 15267
rect 45507 12884 45573 12885
rect 45507 12820 45508 12884
rect 45572 12820 45573 12884
rect 45507 12819 45573 12820
rect 45323 10844 45389 10845
rect 45323 10780 45324 10844
rect 45388 10780 45389 10844
rect 45323 10779 45389 10780
rect 45694 8805 45754 17715
rect 46062 10301 46122 22475
rect 49187 20908 49253 20909
rect 49187 20844 49188 20908
rect 49252 20844 49253 20908
rect 49187 20843 49253 20844
rect 48267 17100 48333 17101
rect 48267 17036 48268 17100
rect 48332 17036 48333 17100
rect 48267 17035 48333 17036
rect 48635 17100 48701 17101
rect 48635 17036 48636 17100
rect 48700 17036 48701 17100
rect 48635 17035 48701 17036
rect 47347 13156 47413 13157
rect 47347 13092 47348 13156
rect 47412 13092 47413 13156
rect 47347 13091 47413 13092
rect 46059 10300 46125 10301
rect 46059 10236 46060 10300
rect 46124 10236 46125 10300
rect 46059 10235 46125 10236
rect 47350 10165 47410 13091
rect 48270 12205 48330 17035
rect 48638 14789 48698 17035
rect 49190 16557 49250 20843
rect 49187 16556 49253 16557
rect 49187 16492 49188 16556
rect 49252 16492 49253 16556
rect 49187 16491 49253 16492
rect 49187 15468 49253 15469
rect 49187 15404 49188 15468
rect 49252 15404 49253 15468
rect 49187 15403 49253 15404
rect 48635 14788 48701 14789
rect 48635 14724 48636 14788
rect 48700 14724 48701 14788
rect 48635 14723 48701 14724
rect 48451 13564 48517 13565
rect 48451 13500 48452 13564
rect 48516 13500 48517 13564
rect 48451 13499 48517 13500
rect 48267 12204 48333 12205
rect 48267 12140 48268 12204
rect 48332 12140 48333 12204
rect 48267 12139 48333 12140
rect 47347 10164 47413 10165
rect 47347 10100 47348 10164
rect 47412 10100 47413 10164
rect 47347 10099 47413 10100
rect 45691 8804 45757 8805
rect 45691 8740 45692 8804
rect 45756 8740 45757 8804
rect 45691 8739 45757 8740
rect 48454 6901 48514 13499
rect 48638 13293 48698 14723
rect 48635 13292 48701 13293
rect 48635 13228 48636 13292
rect 48700 13228 48701 13292
rect 48635 13227 48701 13228
rect 49190 12613 49250 15403
rect 49374 14925 49434 24787
rect 49371 14924 49437 14925
rect 49371 14860 49372 14924
rect 49436 14860 49437 14924
rect 49371 14859 49437 14860
rect 49371 13700 49437 13701
rect 49371 13636 49372 13700
rect 49436 13636 49437 13700
rect 49371 13635 49437 13636
rect 49187 12612 49253 12613
rect 49187 12548 49188 12612
rect 49252 12548 49253 12612
rect 49187 12547 49253 12548
rect 49374 8261 49434 13635
rect 49371 8260 49437 8261
rect 49371 8196 49372 8260
rect 49436 8196 49437 8260
rect 49371 8195 49437 8196
rect 44587 6900 44653 6901
rect 44587 6836 44588 6900
rect 44652 6836 44653 6900
rect 44587 6835 44653 6836
rect 48451 6900 48517 6901
rect 48451 6836 48452 6900
rect 48516 6836 48517 6900
rect 48451 6835 48517 6836
rect 39803 5812 39869 5813
rect 39803 5748 39804 5812
rect 39868 5748 39869 5812
rect 39803 5747 39869 5748
rect 37595 5540 37661 5541
rect 37595 5476 37596 5540
rect 37660 5476 37661 5540
rect 37595 5475 37661 5476
rect 36123 4044 36189 4045
rect 36123 3980 36124 4044
rect 36188 3980 36189 4044
rect 36123 3979 36189 3980
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 49926 2685 49986 27643
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 53419 21316 53485 21317
rect 53419 21252 53420 21316
rect 53484 21252 53485 21316
rect 53419 21251 53485 21252
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 52315 19276 52381 19277
rect 52315 19212 52316 19276
rect 52380 19212 52381 19276
rect 52315 19211 52381 19212
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50843 12884 50909 12885
rect 50843 12820 50844 12884
rect 50908 12820 50909 12884
rect 50843 12819 50909 12820
rect 50846 12450 50906 12819
rect 50846 12390 51274 12450
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 51214 8125 51274 12390
rect 52318 12341 52378 19211
rect 53422 15197 53482 21251
rect 53971 18052 54037 18053
rect 53971 17988 53972 18052
rect 54036 17988 54037 18052
rect 53971 17987 54037 17988
rect 53787 16692 53853 16693
rect 53787 16628 53788 16692
rect 53852 16628 53853 16692
rect 53787 16627 53853 16628
rect 53419 15196 53485 15197
rect 53419 15132 53420 15196
rect 53484 15132 53485 15196
rect 53419 15131 53485 15132
rect 53790 12341 53850 16627
rect 52315 12340 52381 12341
rect 52315 12276 52316 12340
rect 52380 12276 52381 12340
rect 52315 12275 52381 12276
rect 53787 12340 53853 12341
rect 53787 12276 53788 12340
rect 53852 12276 53853 12340
rect 53787 12275 53853 12276
rect 53974 10845 54034 17987
rect 53971 10844 54037 10845
rect 53971 10780 53972 10844
rect 54036 10780 54037 10844
rect 53971 10779 54037 10780
rect 55075 10844 55141 10845
rect 55075 10780 55076 10844
rect 55140 10780 55141 10844
rect 55075 10779 55141 10780
rect 51947 8940 52013 8941
rect 51947 8876 51948 8940
rect 52012 8876 52013 8940
rect 51947 8875 52013 8876
rect 51211 8124 51277 8125
rect 51211 8060 51212 8124
rect 51276 8060 51277 8124
rect 51211 8059 51277 8060
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 51950 5269 52010 8875
rect 55078 6765 55138 10779
rect 55075 6764 55141 6765
rect 55075 6700 55076 6764
rect 55140 6700 55141 6764
rect 55075 6699 55141 6700
rect 51947 5268 52013 5269
rect 51947 5204 51948 5268
rect 52012 5204 52013 5268
rect 51947 5203 52013 5204
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 49923 2684 49989 2685
rect 49923 2620 49924 2684
rect 49988 2620 49989 2684
rect 49923 2619 49989 2620
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 58236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1666464484
transform 1 0 51888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B
timestamp 1666464484
transform 1 0 54280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__C
timestamp 1666464484
transform -1 0 51520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1666464484
transform 1 0 54648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A_N
timestamp 1666464484
transform -1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B
timestamp 1666464484
transform 1 0 57316 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A
timestamp 1666464484
transform 1 0 57132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 1666464484
transform 1 0 56488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1666464484
transform 1 0 52164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A
timestamp 1666464484
transform 1 0 57684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1666464484
transform -1 0 55568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__C
timestamp 1666464484
transform 1 0 57040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A
timestamp 1666464484
transform -1 0 53084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B
timestamp 1666464484
transform 1 0 57408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A2
timestamp 1666464484
transform -1 0 58420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B1
timestamp 1666464484
transform 1 0 57684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__C1
timestamp 1666464484
transform 1 0 56396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A2
timestamp 1666464484
transform 1 0 56856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A3
timestamp 1666464484
transform 1 0 57132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__B1
timestamp 1666464484
transform 1 0 57592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A2
timestamp 1666464484
transform -1 0 57592 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1666464484
transform 1 0 41584 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A
timestamp 1666464484
transform 1 0 42596 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1666464484
transform -1 0 48668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__D_N
timestamp 1666464484
transform 1 0 36708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1666464484
transform 1 0 29072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1666464484
transform 1 0 37996 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1666464484
transform 1 0 41216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B_N
timestamp 1666464484
transform 1 0 40940 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B1
timestamp 1666464484
transform -1 0 38824 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A2
timestamp 1666464484
transform -1 0 32476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B1
timestamp 1666464484
transform 1 0 32844 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__C1
timestamp 1666464484
transform 1 0 32292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A
timestamp 1666464484
transform -1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A0
timestamp 1666464484
transform 1 0 44988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__S
timestamp 1666464484
transform 1 0 44436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__S
timestamp 1666464484
transform 1 0 45172 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A0
timestamp 1666464484
transform 1 0 25392 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__S
timestamp 1666464484
transform 1 0 24840 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A_N
timestamp 1666464484
transform 1 0 43240 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B
timestamp 1666464484
transform 1 0 41400 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A
timestamp 1666464484
transform -1 0 21896 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1666464484
transform 1 0 23736 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1666464484
transform 1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B
timestamp 1666464484
transform -1 0 29256 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A1
timestamp 1666464484
transform 1 0 30544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B
timestamp 1666464484
transform 1 0 33304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A1
timestamp 1666464484
transform 1 0 29532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1666464484
transform -1 0 41952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__B
timestamp 1666464484
transform 1 0 42596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__B
timestamp 1666464484
transform -1 0 29808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A_N
timestamp 1666464484
transform 1 0 28152 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B
timestamp 1666464484
transform 1 0 28060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__B
timestamp 1666464484
transform -1 0 41676 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A2
timestamp 1666464484
transform -1 0 40940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A
timestamp 1666464484
transform 1 0 25852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A2
timestamp 1666464484
transform 1 0 28796 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A
timestamp 1666464484
transform 1 0 26036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B
timestamp 1666464484
transform 1 0 24104 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A2
timestamp 1666464484
transform 1 0 24564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B1_N
timestamp 1666464484
transform 1 0 31740 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1666464484
transform -1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1666464484
transform 1 0 39284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B
timestamp 1666464484
transform 1 0 40020 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__B
timestamp 1666464484
transform 1 0 32936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__B1
timestamp 1666464484
transform -1 0 41216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__C1
timestamp 1666464484
transform 1 0 40664 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A
timestamp 1666464484
transform -1 0 23828 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A
timestamp 1666464484
transform 1 0 34500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__C
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__C1
timestamp 1666464484
transform 1 0 27876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__A
timestamp 1666464484
transform -1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__B
timestamp 1666464484
transform 1 0 41032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1666464484
transform 1 0 39100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A1
timestamp 1666464484
transform 1 0 28244 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A1
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1666464484
transform 1 0 27876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A_N
timestamp 1666464484
transform 1 0 29072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__B
timestamp 1666464484
transform -1 0 36892 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__B1
timestamp 1666464484
transform 1 0 28520 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A1_N
timestamp 1666464484
transform -1 0 27416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A1
timestamp 1666464484
transform -1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B2
timestamp 1666464484
transform -1 0 24564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1666464484
transform 1 0 30636 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A1
timestamp 1666464484
transform 1 0 29716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1666464484
transform -1 0 44620 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A3
timestamp 1666464484
transform 1 0 26956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__B1
timestamp 1666464484
transform 1 0 25944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1666464484
transform 1 0 26128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A1_N
timestamp 1666464484
transform 1 0 26680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A2_N
timestamp 1666464484
transform -1 0 25484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__C1
timestamp 1666464484
transform -1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1666464484
transform 1 0 28612 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__B1
timestamp 1666464484
transform 1 0 29900 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1666464484
transform 1 0 28612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__B
timestamp 1666464484
transform 1 0 29164 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A
timestamp 1666464484
transform 1 0 31096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A0
timestamp 1666464484
transform -1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__S1
timestamp 1666464484
transform -1 0 27324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A1
timestamp 1666464484
transform -1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__B1
timestamp 1666464484
transform 1 0 23920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A1_N
timestamp 1666464484
transform -1 0 24012 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A2
timestamp 1666464484
transform 1 0 31648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A1
timestamp 1666464484
transform 1 0 29072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A
timestamp 1666464484
transform -1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A
timestamp 1666464484
transform 1 0 27140 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__B
timestamp 1666464484
transform 1 0 29072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A1
timestamp 1666464484
transform 1 0 26864 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B
timestamp 1666464484
transform 1 0 34224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A
timestamp 1666464484
transform 1 0 24104 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A1
timestamp 1666464484
transform 1 0 25116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__B1
timestamp 1666464484
transform -1 0 24380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__A1
timestamp 1666464484
transform 1 0 25668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A2
timestamp 1666464484
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__B1
timestamp 1666464484
transform 1 0 26312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__B1
timestamp 1666464484
transform -1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A1
timestamp 1666464484
transform 1 0 26496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__B1
timestamp 1666464484
transform 1 0 30544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A
timestamp 1666464484
transform -1 0 29900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__A1
timestamp 1666464484
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B
timestamp 1666464484
transform 1 0 34224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A1
timestamp 1666464484
transform 1 0 36800 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B2
timestamp 1666464484
transform 1 0 36156 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B
timestamp 1666464484
transform 1 0 31648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B
timestamp 1666464484
transform 1 0 33304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A2
timestamp 1666464484
transform -1 0 33304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B1
timestamp 1666464484
transform 1 0 32568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__B
timestamp 1666464484
transform -1 0 38824 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A
timestamp 1666464484
transform 1 0 39192 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A1
timestamp 1666464484
transform 1 0 31740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A
timestamp 1666464484
transform 1 0 28520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1666464484
transform -1 0 58236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__A
timestamp 1666464484
transform 1 0 33948 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__B
timestamp 1666464484
transform -1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__B
timestamp 1666464484
transform 1 0 41400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A1
timestamp 1666464484
transform 1 0 35420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A1
timestamp 1666464484
transform 1 0 33396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A1_N
timestamp 1666464484
transform 1 0 33120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A2_N
timestamp 1666464484
transform 1 0 35972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B1
timestamp 1666464484
transform -1 0 36708 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B2
timestamp 1666464484
transform 1 0 34868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1666464484
transform 1 0 34224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__B1
timestamp 1666464484
transform 1 0 34868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1666464484
transform 1 0 33028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A
timestamp 1666464484
transform -1 0 36248 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__A1
timestamp 1666464484
transform 1 0 40848 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1666464484
transform -1 0 41400 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__B
timestamp 1666464484
transform 1 0 40940 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__B
timestamp 1666464484
transform 1 0 40296 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__S
timestamp 1666464484
transform 1 0 41584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A
timestamp 1666464484
transform -1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A1
timestamp 1666464484
transform 1 0 37444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__B2
timestamp 1666464484
transform 1 0 37076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 1666464484
transform 1 0 40480 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__A
timestamp 1666464484
transform 1 0 36800 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A1
timestamp 1666464484
transform 1 0 39284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__B1
timestamp 1666464484
transform 1 0 35420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A
timestamp 1666464484
transform 1 0 34316 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__A
timestamp 1666464484
transform -1 0 37904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 1666464484
transform 1 0 39284 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__A_N
timestamp 1666464484
transform -1 0 42320 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__C
timestamp 1666464484
transform 1 0 38916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__A2
timestamp 1666464484
transform 1 0 35972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A
timestamp 1666464484
transform 1 0 35972 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__C
timestamp 1666464484
transform 1 0 38272 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__B1
timestamp 1666464484
transform -1 0 38824 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__B1
timestamp 1666464484
transform -1 0 40112 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__B2
timestamp 1666464484
transform -1 0 39376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A0
timestamp 1666464484
transform 1 0 40020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__A2
timestamp 1666464484
transform 1 0 37444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__A
timestamp 1666464484
transform 1 0 36340 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__A
timestamp 1666464484
transform -1 0 41952 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A
timestamp 1666464484
transform 1 0 56580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A
timestamp 1666464484
transform 1 0 45724 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__A
timestamp 1666464484
transform 1 0 53452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__A
timestamp 1666464484
transform 1 0 42320 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__A
timestamp 1666464484
transform 1 0 50324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__A
timestamp 1666464484
transform 1 0 56028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__A
timestamp 1666464484
transform 1 0 45172 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__A
timestamp 1666464484
transform 1 0 51612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__A1
timestamp 1666464484
transform 1 0 45816 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__B
timestamp 1666464484
transform 1 0 56488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__A
timestamp 1666464484
transform 1 0 56856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__A
timestamp 1666464484
transform 1 0 55936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__A2
timestamp 1666464484
transform -1 0 56948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__B2
timestamp 1666464484
transform 1 0 50140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1522__A1
timestamp 1666464484
transform 1 0 49496 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__A
timestamp 1666464484
transform 1 0 53544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1527__A
timestamp 1666464484
transform 1 0 47748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1527__B
timestamp 1666464484
transform 1 0 45908 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1529__A1
timestamp 1666464484
transform -1 0 54188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1530__A2
timestamp 1666464484
transform 1 0 50600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1532__A2
timestamp 1666464484
transform 1 0 48852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1532__A3
timestamp 1666464484
transform 1 0 51244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1533__A
timestamp 1666464484
transform 1 0 42688 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__A
timestamp 1666464484
transform 1 0 47472 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__A
timestamp 1666464484
transform 1 0 43240 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1536__A1
timestamp 1666464484
transform 1 0 48760 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__A_N
timestamp 1666464484
transform -1 0 51244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__A
timestamp 1666464484
transform 1 0 57224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__A2
timestamp 1666464484
transform 1 0 45172 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1543__A1
timestamp 1666464484
transform 1 0 48300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1545__A
timestamp 1666464484
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1547__A
timestamp 1666464484
transform -1 0 48760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1548__A
timestamp 1666464484
transform -1 0 49312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1549__B1
timestamp 1666464484
transform 1 0 54096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1552__A
timestamp 1666464484
transform 1 0 54740 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__A
timestamp 1666464484
transform -1 0 53084 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__B
timestamp 1666464484
transform 1 0 53452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1557__A1
timestamp 1666464484
transform 1 0 54740 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__A
timestamp 1666464484
transform -1 0 42044 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__A1
timestamp 1666464484
transform 1 0 53728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1560__B2
timestamp 1666464484
transform 1 0 52716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1561__A
timestamp 1666464484
transform 1 0 46460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__A_N
timestamp 1666464484
transform 1 0 48852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__B
timestamp 1666464484
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1577__A1
timestamp 1666464484
transform -1 0 52348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__A
timestamp 1666464484
transform 1 0 51520 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__A2
timestamp 1666464484
transform 1 0 47380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1581__B
timestamp 1666464484
transform -1 0 46828 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1584__B
timestamp 1666464484
transform -1 0 57132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1586__B1
timestamp 1666464484
transform -1 0 50784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1588__A2
timestamp 1666464484
transform 1 0 55384 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1589__B
timestamp 1666464484
transform 1 0 54832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1591__B1
timestamp 1666464484
transform 1 0 51152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1597__C
timestamp 1666464484
transform 1 0 47748 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1598__B1
timestamp 1666464484
transform -1 0 47196 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__A2
timestamp 1666464484
transform 1 0 49588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__B1
timestamp 1666464484
transform 1 0 53820 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1602__A
timestamp 1666464484
transform 1 0 46552 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1603__B1
timestamp 1666464484
transform 1 0 47748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__A
timestamp 1666464484
transform 1 0 46368 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__B1
timestamp 1666464484
transform 1 0 48944 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__A1
timestamp 1666464484
transform 1 0 56304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1620__B
timestamp 1666464484
transform 1 0 44068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1622__A
timestamp 1666464484
transform 1 0 46644 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1627__A
timestamp 1666464484
transform -1 0 57960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1630__A1
timestamp 1666464484
transform 1 0 47104 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1630__B1
timestamp 1666464484
transform 1 0 49496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1634__B1
timestamp 1666464484
transform 1 0 47472 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1635__A1
timestamp 1666464484
transform 1 0 43240 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1636__A1
timestamp 1666464484
transform 1 0 51244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1636__B1
timestamp 1666464484
transform 1 0 52256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1637__B_N
timestamp 1666464484
transform 1 0 46276 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1639__B
timestamp 1666464484
transform 1 0 49036 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1640__B
timestamp 1666464484
transform 1 0 45724 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1649__B1
timestamp 1666464484
transform -1 0 47288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1650__C
timestamp 1666464484
transform 1 0 45816 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1656__A
timestamp 1666464484
transform -1 0 44528 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1667__B
timestamp 1666464484
transform 1 0 46184 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1667__C
timestamp 1666464484
transform -1 0 48484 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1668__A1
timestamp 1666464484
transform 1 0 49588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1669__B1
timestamp 1666464484
transform -1 0 48484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1670__A2
timestamp 1666464484
transform 1 0 50048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1671__A1
timestamp 1666464484
transform -1 0 48484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1673__A1
timestamp 1666464484
transform 1 0 42872 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1673__A2
timestamp 1666464484
transform 1 0 44988 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1673__B1
timestamp 1666464484
transform 1 0 43424 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1679__A
timestamp 1666464484
transform 1 0 46276 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1681__A1
timestamp 1666464484
transform 1 0 44436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1682__A1
timestamp 1666464484
transform 1 0 42412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1685__A1
timestamp 1666464484
transform 1 0 52164 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1693__A1
timestamp 1666464484
transform 1 0 57040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1693__B1
timestamp 1666464484
transform -1 0 54372 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1693__B2
timestamp 1666464484
transform -1 0 54004 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1693__C1
timestamp 1666464484
transform -1 0 55568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1695__A
timestamp 1666464484
transform -1 0 58328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1695__B
timestamp 1666464484
transform -1 0 58236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1696__B2
timestamp 1666464484
transform 1 0 56672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1697__A
timestamp 1666464484
transform 1 0 55476 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1698__A1
timestamp 1666464484
transform 1 0 56948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1699__A1_N
timestamp 1666464484
transform 1 0 56396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1702__A
timestamp 1666464484
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1712__A2
timestamp 1666464484
transform 1 0 46552 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1712__A3
timestamp 1666464484
transform 1 0 47104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1713__A1
timestamp 1666464484
transform 1 0 45172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1713__A2
timestamp 1666464484
transform 1 0 42596 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1715__A1
timestamp 1666464484
transform 1 0 49680 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1716__A2
timestamp 1666464484
transform 1 0 44344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1721__A
timestamp 1666464484
transform 1 0 55752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1721__B
timestamp 1666464484
transform 1 0 56304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1723__A
timestamp 1666464484
transform 1 0 55476 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1723__B
timestamp 1666464484
transform 1 0 56028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1724__A
timestamp 1666464484
transform -1 0 56764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1726__A
timestamp 1666464484
transform 1 0 57132 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1727__A1
timestamp 1666464484
transform 1 0 54372 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1727__C1
timestamp 1666464484
transform 1 0 55016 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1733__A1
timestamp 1666464484
transform -1 0 49128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1734__B1
timestamp 1666464484
transform 1 0 54832 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1743__A1
timestamp 1666464484
transform 1 0 55016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1743__A2
timestamp 1666464484
transform 1 0 54832 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1743__A3
timestamp 1666464484
transform -1 0 54464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1743__C1
timestamp 1666464484
transform 1 0 56948 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1744__A1
timestamp 1666464484
transform 1 0 56120 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1744__B1
timestamp 1666464484
transform 1 0 56672 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1745__A
timestamp 1666464484
transform 1 0 42780 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1746__A
timestamp 1666464484
transform 1 0 49588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1747__B
timestamp 1666464484
transform 1 0 47748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1748__A
timestamp 1666464484
transform 1 0 44068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1749__A1
timestamp 1666464484
transform 1 0 54832 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1751__B1
timestamp 1666464484
transform 1 0 49588 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1762__A
timestamp 1666464484
transform 1 0 46920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1766__B
timestamp 1666464484
transform 1 0 51520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1766__C_N
timestamp 1666464484
transform 1 0 52900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1767__A1
timestamp 1666464484
transform 1 0 52164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1767__C1
timestamp 1666464484
transform 1 0 51244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1768__A
timestamp 1666464484
transform 1 0 50784 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1768__B
timestamp 1666464484
transform 1 0 51888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1769__A1
timestamp 1666464484
transform -1 0 51520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1770__A1
timestamp 1666464484
transform -1 0 48208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1781__A
timestamp 1666464484
transform 1 0 50324 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1782__A
timestamp 1666464484
transform 1 0 56212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1783__A2
timestamp 1666464484
transform -1 0 58236 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1785__A
timestamp 1666464484
transform 1 0 57316 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1786__A1
timestamp 1666464484
transform 1 0 50692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1787__A
timestamp 1666464484
transform 1 0 57040 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1788__A1
timestamp 1666464484
transform 1 0 56764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1798__A1
timestamp 1666464484
transform 1 0 55936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1799__A1
timestamp 1666464484
transform 1 0 57960 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1800__A
timestamp 1666464484
transform -1 0 57040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1803__A1
timestamp 1666464484
transform 1 0 54372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1803__B2
timestamp 1666464484
transform -1 0 54004 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1808__A1
timestamp 1666464484
transform 1 0 42688 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1809__A
timestamp 1666464484
transform 1 0 41952 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1810__A1
timestamp 1666464484
transform -1 0 42872 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1810__A2
timestamp 1666464484
transform 1 0 45264 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1811__B2
timestamp 1666464484
transform 1 0 46828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1817__A
timestamp 1666464484
transform 1 0 57040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1818__A1
timestamp 1666464484
transform 1 0 57776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1820__A1
timestamp 1666464484
transform 1 0 56580 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1829__A
timestamp 1666464484
transform -1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1830__A1
timestamp 1666464484
transform 1 0 56856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1831__A1
timestamp 1666464484
transform -1 0 58236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1831__A2
timestamp 1666464484
transform -1 0 58236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1831__B1
timestamp 1666464484
transform 1 0 57500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1833__A1
timestamp 1666464484
transform -1 0 58236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1836__A
timestamp 1666464484
transform -1 0 56580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1836__B
timestamp 1666464484
transform 1 0 53728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1838__A
timestamp 1666464484
transform 1 0 56028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1839__A
timestamp 1666464484
transform 1 0 56580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1840__A
timestamp 1666464484
transform -1 0 58236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1842__A3
timestamp 1666464484
transform 1 0 56580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1848__A1
timestamp 1666464484
transform 1 0 57408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1848__A3
timestamp 1666464484
transform 1 0 55936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1862__B
timestamp 1666464484
transform 1 0 56948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1864__A1
timestamp 1666464484
transform 1 0 57224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1864__A2
timestamp 1666464484
transform -1 0 57684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1864__A3
timestamp 1666464484
transform -1 0 58236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1865__A
timestamp 1666464484
transform -1 0 58236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1872__A2
timestamp 1666464484
transform 1 0 57224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1873__A
timestamp 1666464484
transform -1 0 56856 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1873__B
timestamp 1666464484
transform 1 0 57224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1873__C
timestamp 1666464484
transform 1 0 56488 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1878__A1
timestamp 1666464484
transform 1 0 52900 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1878__B2
timestamp 1666464484
transform -1 0 49864 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1878__C1
timestamp 1666464484
transform 1 0 55292 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1880__A2
timestamp 1666464484
transform -1 0 57408 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1882__S
timestamp 1666464484
transform 1 0 56580 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1892__A1
timestamp 1666464484
transform 1 0 57132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1892__A2
timestamp 1666464484
transform -1 0 58236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1893__B1
timestamp 1666464484
transform 1 0 57776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1894__A
timestamp 1666464484
transform -1 0 58236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1895__A1
timestamp 1666464484
transform -1 0 54556 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1898__B1
timestamp 1666464484
transform -1 0 57316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1907__A0
timestamp 1666464484
transform 1 0 57776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1919__A1
timestamp 1666464484
transform -1 0 52256 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1919__A2
timestamp 1666464484
transform -1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1920__B2
timestamp 1666464484
transform 1 0 56856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1927__A1
timestamp 1666464484
transform -1 0 58236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1938__A1
timestamp 1666464484
transform 1 0 54648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1958__A0
timestamp 1666464484
transform -1 0 50232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1958__S
timestamp 1666464484
transform -1 0 55660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1960__A1
timestamp 1666464484
transform 1 0 45632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1960__S
timestamp 1666464484
transform 1 0 45172 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1963__A0
timestamp 1666464484
transform -1 0 47932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1963__S
timestamp 1666464484
transform -1 0 46552 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1965__B
timestamp 1666464484
transform 1 0 46092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1966__A
timestamp 1666464484
transform 1 0 44252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1966__B
timestamp 1666464484
transform 1 0 45172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1967__A
timestamp 1666464484
transform 1 0 41952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1968__A1_N
timestamp 1666464484
transform 1 0 46276 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1968__B1
timestamp 1666464484
transform -1 0 44344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1969__A1
timestamp 1666464484
transform 1 0 45724 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1969__A3
timestamp 1666464484
transform 1 0 47104 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1969__B1
timestamp 1666464484
transform 1 0 46184 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1972__A
timestamp 1666464484
transform 1 0 49220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1973__A1
timestamp 1666464484
transform -1 0 49220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1973__B1
timestamp 1666464484
transform -1 0 48208 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1974__A
timestamp 1666464484
transform -1 0 47012 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1974__B
timestamp 1666464484
transform 1 0 47748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1975__A1
timestamp 1666464484
transform -1 0 50416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1975__A2
timestamp 1666464484
transform 1 0 50784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1976__A1
timestamp 1666464484
transform -1 0 45448 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1976__B2
timestamp 1666464484
transform 1 0 51428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1977__A1
timestamp 1666464484
transform -1 0 49680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1978__B
timestamp 1666464484
transform 1 0 45080 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1982__A1
timestamp 1666464484
transform -1 0 41768 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1986__A2
timestamp 1666464484
transform 1 0 41860 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1986__B1
timestamp 1666464484
transform 1 0 42044 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1990__A
timestamp 1666464484
transform -1 0 21620 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1991__A
timestamp 1666464484
transform -1 0 55292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1991__B
timestamp 1666464484
transform -1 0 55660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1992__A1
timestamp 1666464484
transform -1 0 49036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2011__RESET_B
timestamp 1666464484
transform 1 0 24564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2012__D
timestamp 1666464484
transform 1 0 23184 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2012__RESET_B
timestamp 1666464484
transform 1 0 25576 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2013__CLK
timestamp 1666464484
transform 1 0 46828 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2013__RESET_B
timestamp 1666464484
transform 1 0 45172 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2015__CLK
timestamp 1666464484
transform 1 0 45724 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2015__RESET_B
timestamp 1666464484
transform 1 0 42688 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2017__D
timestamp 1666464484
transform 1 0 23828 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2017__RESET_B
timestamp 1666464484
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2019__RESET_B
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2020__CLK
timestamp 1666464484
transform 1 0 43516 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2020__RESET_B
timestamp 1666464484
transform -1 0 41768 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2021__CLK
timestamp 1666464484
transform 1 0 44804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2021__RESET_B
timestamp 1666464484
transform 1 0 41952 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_CLK_A
timestamp 1666464484
transform -1 0 48116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout42_A
timestamp 1666464484
transform -1 0 54740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout43_A
timestamp 1666464484
transform 1 0 42136 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout45_A
timestamp 1666464484
transform -1 0 46000 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout46_A
timestamp 1666464484
transform 1 0 41308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout47_A
timestamp 1666464484
transform -1 0 47932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout48_A
timestamp 1666464484
transform -1 0 37628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout49_A
timestamp 1666464484
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 31832 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output4_A
timestamp 1666464484
transform -1 0 2484 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_A
timestamp 1666464484
transform 1 0 56856 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output6_A
timestamp 1666464484
transform -1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output8_A
timestamp 1666464484
transform 1 0 4692 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output9_A
timestamp 1666464484
transform -1 0 2484 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output10_A
timestamp 1666464484
transform -1 0 49588 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_A
timestamp 1666464484
transform -1 0 57684 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output14_A
timestamp 1666464484
transform 1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output15_A
timestamp 1666464484
transform 1 0 2300 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output16_A
timestamp 1666464484
transform -1 0 2484 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output17_A
timestamp 1666464484
transform 1 0 37536 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output19_A
timestamp 1666464484
transform 1 0 2300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output20_A
timestamp 1666464484
transform 1 0 57408 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output21_A
timestamp 1666464484
transform 1 0 15916 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_A
timestamp 1666464484
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output23_A
timestamp 1666464484
transform -1 0 2484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output25_A
timestamp 1666464484
transform 1 0 10488 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output26_A
timestamp 1666464484
transform 1 0 2300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_A
timestamp 1666464484
transform -1 0 54188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_A
timestamp 1666464484
transform -1 0 44160 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output29_A
timestamp 1666464484
transform -1 0 58236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 1666464484
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1666464484
transform 1 0 22724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output32_A
timestamp 1666464484
transform -1 0 58236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output33_A
timestamp 1666464484
transform 1 0 28520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output34_A
timestamp 1666464484
transform -1 0 57684 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output35_A
timestamp 1666464484
transform 1 0 57408 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output36_A
timestamp 1666464484
transform 1 0 22724 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output37_A
timestamp 1666464484
transform 1 0 27876 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output39_A
timestamp 1666464484
transform 1 0 2300 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output40_A
timestamp 1666464484
transform 1 0 2300 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1666464484
transform -1 0 56856 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61
timestamp 1666464484
transform 1 0 6716 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7820 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1666464484
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1666464484
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1666464484
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1666464484
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1666464484
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1666464484
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1666464484
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1666464484
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1666464484
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1666464484
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1666464484
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1666464484
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1666464484
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_231
timestamp 1666464484
transform 1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1666464484
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1666464484
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1666464484
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1666464484
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_289
timestamp 1666464484
transform 1 0 27692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_294
timestamp 1666464484
transform 1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_300
timestamp 1666464484
transform 1 0 28704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1666464484
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_313
timestamp 1666464484
transform 1 0 29900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_318
timestamp 1666464484
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_328
timestamp 1666464484
transform 1 0 31280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1666464484
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_343 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1666464484
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1666464484
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_383
timestamp 1666464484
transform 1 0 36340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1666464484
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1666464484
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_427
timestamp 1666464484
transform 1 0 40388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_433
timestamp 1666464484
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_439
timestamp 1666464484
transform 1 0 41492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1666464484
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 1666464484
transform 1 0 44436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1666464484
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_477
timestamp 1666464484
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_482
timestamp 1666464484
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_488
timestamp 1666464484
transform 1 0 46000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1666464484
transform 1 0 46552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1666464484
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_509
timestamp 1666464484
transform 1 0 47932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1666464484
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_521
timestamp 1666464484
transform 1 0 49036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_527
timestamp 1666464484
transform 1 0 49588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1666464484
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1666464484
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1666464484
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_545
timestamp 1666464484
transform 1 0 51244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_551
timestamp 1666464484
transform 1 0 51796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1666464484
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_565
timestamp 1666464484
transform 1 0 53084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1666464484
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_577
timestamp 1666464484
transform 1 0 54188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1666464484
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_597
timestamp 1666464484
transform 1 0 56028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_602
timestamp 1666464484
transform 1 0 56488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_608
timestamp 1666464484
transform 1 0 57040 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1666464484
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1666464484
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1666464484
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1666464484
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1666464484
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1666464484
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1666464484
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1666464484
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1666464484
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1666464484
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1666464484
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1666464484
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1666464484
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1666464484
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1666464484
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1666464484
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1666464484
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_301
timestamp 1666464484
transform 1 0 28796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1666464484
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_312
timestamp 1666464484
transform 1 0 29808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_321
timestamp 1666464484
transform 1 0 30636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1666464484
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666464484
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_348
timestamp 1666464484
transform 1 0 33120 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_376
timestamp 1666464484
transform 1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1666464484
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_397
timestamp 1666464484
transform 1 0 37628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_403
timestamp 1666464484
transform 1 0 38180 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_432
timestamp 1666464484
transform 1 0 40848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_436
timestamp 1666464484
transform 1 0 41216 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1666464484
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666464484
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_474
timestamp 1666464484
transform 1 0 44712 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_501
timestamp 1666464484
transform 1 0 47196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666464484
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_509
timestamp 1666464484
transform 1 0 47932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1666464484
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_521
timestamp 1666464484
transform 1 0 49036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_527
timestamp 1666464484
transform 1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_531
timestamp 1666464484
transform 1 0 49956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_534
timestamp 1666464484
transform 1 0 50232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_540
timestamp 1666464484
transform 1 0 50784 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_548
timestamp 1666464484
transform 1 0 51520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_554
timestamp 1666464484
transform 1 0 52072 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_565
timestamp 1666464484
transform 1 0 53084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1666464484
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_577
timestamp 1666464484
transform 1 0 54188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_583
timestamp 1666464484
transform 1 0 54740 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_589
timestamp 1666464484
transform 1 0 55292 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_601
timestamp 1666464484
transform 1 0 56396 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_613
timestamp 1666464484
transform 1 0 57500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_617
timestamp 1666464484
transform 1 0 57868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1666464484
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1666464484
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1666464484
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1666464484
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1666464484
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1666464484
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1666464484
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1666464484
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1666464484
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1666464484
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1666464484
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1666464484
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1666464484
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1666464484
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1666464484
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1666464484
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1666464484
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_289
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_297
timestamp 1666464484
transform 1 0 28428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1666464484
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_319
timestamp 1666464484
transform 1 0 30452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_329
timestamp 1666464484
transform 1 0 31372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_335
timestamp 1666464484
transform 1 0 31924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_346
timestamp 1666464484
transform 1 0 32936 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_352
timestamp 1666464484
transform 1 0 33488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1666464484
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_371
timestamp 1666464484
transform 1 0 35236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1666464484
transform 1 0 37720 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_409
timestamp 1666464484
transform 1 0 38732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1666464484
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1666464484
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_425
timestamp 1666464484
transform 1 0 40204 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1666464484
transform 1 0 40572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_456
timestamp 1666464484
transform 1 0 43056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_464
timestamp 1666464484
transform 1 0 43792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1666464484
transform 1 0 44344 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666464484
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_481
timestamp 1666464484
transform 1 0 45356 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_485
timestamp 1666464484
transform 1 0 45724 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_506
timestamp 1666464484
transform 1 0 47656 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_512
timestamp 1666464484
transform 1 0 48208 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_518
timestamp 1666464484
transform 1 0 48760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1666464484
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1666464484
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_537
timestamp 1666464484
transform 1 0 50508 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_543
timestamp 1666464484
transform 1 0 51060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_566
timestamp 1666464484
transform 1 0 53176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_572
timestamp 1666464484
transform 1 0 53728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_578
timestamp 1666464484
transform 1 0 54280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_584
timestamp 1666464484
transform 1 0 54832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_589
timestamp 1666464484
transform 1 0 55292 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_593
timestamp 1666464484
transform 1 0 55660 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_605
timestamp 1666464484
transform 1 0 56764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_617
timestamp 1666464484
transform 1 0 57868 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1666464484
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1666464484
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1666464484
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1666464484
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1666464484
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1666464484
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1666464484
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1666464484
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1666464484
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1666464484
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1666464484
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1666464484
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1666464484
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1666464484
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_289
timestamp 1666464484
transform 1 0 27692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_299
timestamp 1666464484
transform 1 0 28612 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_303
timestamp 1666464484
transform 1 0 28980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_306
timestamp 1666464484
transform 1 0 29256 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_317
timestamp 1666464484
transform 1 0 30268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_323
timestamp 1666464484
transform 1 0 30820 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_327
timestamp 1666464484
transform 1 0 31188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1666464484
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_346
timestamp 1666464484
transform 1 0 32936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_352
timestamp 1666464484
transform 1 0 33488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_363
timestamp 1666464484
transform 1 0 34500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_390
timestamp 1666464484
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_416
timestamp 1666464484
transform 1 0 39376 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_440
timestamp 1666464484
transform 1 0 41584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_446
timestamp 1666464484
transform 1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_453
timestamp 1666464484
transform 1 0 42780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_457
timestamp 1666464484
transform 1 0 43148 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_481
timestamp 1666464484
transform 1 0 45356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_487
timestamp 1666464484
transform 1 0 45908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_493
timestamp 1666464484
transform 1 0 46460 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1666464484
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_516
timestamp 1666464484
transform 1 0 48576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_522
timestamp 1666464484
transform 1 0 49128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_528
timestamp 1666464484
transform 1 0 49680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_534
timestamp 1666464484
transform 1 0 50232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_540
timestamp 1666464484
transform 1 0 50784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_546
timestamp 1666464484
transform 1 0 51336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_554
timestamp 1666464484
transform 1 0 52072 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_557
timestamp 1666464484
transform 1 0 52348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_561
timestamp 1666464484
transform 1 0 52716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_568
timestamp 1666464484
transform 1 0 53360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_574
timestamp 1666464484
transform 1 0 53912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_580
timestamp 1666464484
transform 1 0 54464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_586
timestamp 1666464484
transform 1 0 55016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_592
timestamp 1666464484
transform 1 0 55568 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_598
timestamp 1666464484
transform 1 0 56120 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_610
timestamp 1666464484
transform 1 0 57224 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1666464484
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1666464484
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1666464484
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1666464484
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1666464484
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1666464484
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1666464484
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1666464484
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_265
timestamp 1666464484
transform 1 0 25484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_271
timestamp 1666464484
transform 1 0 26036 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_274
timestamp 1666464484
transform 1 0 26312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_280
timestamp 1666464484
transform 1 0 26864 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_286
timestamp 1666464484
transform 1 0 27416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_298
timestamp 1666464484
transform 1 0 28520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_302
timestamp 1666464484
transform 1 0 28888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666464484
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_317
timestamp 1666464484
transform 1 0 30268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_329
timestamp 1666464484
transform 1 0 31372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_335
timestamp 1666464484
transform 1 0 31924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_346
timestamp 1666464484
transform 1 0 32936 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_354
timestamp 1666464484
transform 1 0 33672 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1666464484
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_373
timestamp 1666464484
transform 1 0 35420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_400
timestamp 1666464484
transform 1 0 37904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_408
timestamp 1666464484
transform 1 0 38640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_415
timestamp 1666464484
transform 1 0 39284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666464484
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_421
timestamp 1666464484
transform 1 0 39836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_445
timestamp 1666464484
transform 1 0 42044 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_455
timestamp 1666464484
transform 1 0 42964 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_465
timestamp 1666464484
transform 1 0 43884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_471
timestamp 1666464484
transform 1 0 44436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666464484
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1666464484
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_481
timestamp 1666464484
transform 1 0 45356 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_487
timestamp 1666464484
transform 1 0 45908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_493
timestamp 1666464484
transform 1 0 46460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_499
timestamp 1666464484
transform 1 0 47012 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1666464484
transform 1 0 47564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_511
timestamp 1666464484
transform 1 0 48116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_517
timestamp 1666464484
transform 1 0 48668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_523
timestamp 1666464484
transform 1 0 49220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 1666464484
transform 1 0 49772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_533
timestamp 1666464484
transform 1 0 50140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_544
timestamp 1666464484
transform 1 0 51152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_550
timestamp 1666464484
transform 1 0 51704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_556
timestamp 1666464484
transform 1 0 52256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_563
timestamp 1666464484
transform 1 0 52900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_573
timestamp 1666464484
transform 1 0 53820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_579
timestamp 1666464484
transform 1 0 54372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_585
timestamp 1666464484
transform 1 0 54924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_589
timestamp 1666464484
transform 1 0 55292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_593
timestamp 1666464484
transform 1 0 55660 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_599
timestamp 1666464484
transform 1 0 56212 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_605
timestamp 1666464484
transform 1 0 56764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_617
timestamp 1666464484
transform 1 0 57868 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1666464484
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1666464484
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1666464484
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1666464484
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1666464484
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1666464484
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_261
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_269
timestamp 1666464484
transform 1 0 25852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1666464484
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_291
timestamp 1666464484
transform 1 0 27876 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_299
timestamp 1666464484
transform 1 0 28612 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_305
timestamp 1666464484
transform 1 0 29164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1666464484
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_322
timestamp 1666464484
transform 1 0 30728 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_334
timestamp 1666464484
transform 1 0 31832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_350
timestamp 1666464484
transform 1 0 33304 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_357
timestamp 1666464484
transform 1 0 33948 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_383
timestamp 1666464484
transform 1 0 36340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_389
timestamp 1666464484
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1666464484
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_430
timestamp 1666464484
transform 1 0 40664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1666464484
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666464484
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_474
timestamp 1666464484
transform 1 0 44712 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_480
timestamp 1666464484
transform 1 0 45264 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_486
timestamp 1666464484
transform 1 0 45816 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_492
timestamp 1666464484
transform 1 0 46368 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_496
timestamp 1666464484
transform 1 0 46736 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1666464484
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_509
timestamp 1666464484
transform 1 0 47932 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_520
timestamp 1666464484
transform 1 0 48944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_530
timestamp 1666464484
transform 1 0 49864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_536
timestamp 1666464484
transform 1 0 50416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_542
timestamp 1666464484
transform 1 0 50968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_550
timestamp 1666464484
transform 1 0 51704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_558
timestamp 1666464484
transform 1 0 52440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_561
timestamp 1666464484
transform 1 0 52716 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_569
timestamp 1666464484
transform 1 0 53452 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_575
timestamp 1666464484
transform 1 0 54004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_579
timestamp 1666464484
transform 1 0 54372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_586
timestamp 1666464484
transform 1 0 55016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_592
timestamp 1666464484
transform 1 0 55568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_598
timestamp 1666464484
transform 1 0 56120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_604
timestamp 1666464484
transform 1 0 56672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_610
timestamp 1666464484
transform 1 0 57224 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1666464484
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_9
timestamp 1666464484
transform 1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1666464484
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1666464484
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1666464484
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1666464484
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_261
timestamp 1666464484
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_265
timestamp 1666464484
transform 1 0 25484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_277
timestamp 1666464484
transform 1 0 26588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_291
timestamp 1666464484
transform 1 0 27876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1666464484
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1666464484
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_319
timestamp 1666464484
transform 1 0 30452 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_327
timestamp 1666464484
transform 1 0 31188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_336
timestamp 1666464484
transform 1 0 32016 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_344
timestamp 1666464484
transform 1 0 32752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_353
timestamp 1666464484
transform 1 0 33580 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_359
timestamp 1666464484
transform 1 0 34132 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_372
timestamp 1666464484
transform 1 0 35328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_384
timestamp 1666464484
transform 1 0 36432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_397
timestamp 1666464484
transform 1 0 37628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_409
timestamp 1666464484
transform 1 0 38732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_416
timestamp 1666464484
transform 1 0 39376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_425
timestamp 1666464484
transform 1 0 40204 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_433
timestamp 1666464484
transform 1 0 40940 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_442
timestamp 1666464484
transform 1 0 41768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_448
timestamp 1666464484
transform 1 0 42320 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_461
timestamp 1666464484
transform 1 0 43516 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_465
timestamp 1666464484
transform 1 0 43884 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_470
timestamp 1666464484
transform 1 0 44344 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_477
timestamp 1666464484
transform 1 0 44988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_485
timestamp 1666464484
transform 1 0 45724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_491
timestamp 1666464484
transform 1 0 46276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_495
timestamp 1666464484
transform 1 0 46644 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_504
timestamp 1666464484
transform 1 0 47472 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_519
timestamp 1666464484
transform 1 0 48852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_533
timestamp 1666464484
transform 1 0 50140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_543
timestamp 1666464484
transform 1 0 51060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_549
timestamp 1666464484
transform 1 0 51612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_559
timestamp 1666464484
transform 1 0 52532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_569
timestamp 1666464484
transform 1 0 53452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_586
timestamp 1666464484
transform 1 0 55016 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_589
timestamp 1666464484
transform 1 0 55292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_593
timestamp 1666464484
transform 1 0 55660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_599
timestamp 1666464484
transform 1 0 56212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_605
timestamp 1666464484
transform 1 0 56764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_611
timestamp 1666464484
transform 1 0 57316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_617
timestamp 1666464484
transform 1 0 57868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_623
timestamp 1666464484
transform 1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1666464484
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1666464484
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1666464484
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1666464484
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1666464484
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1666464484
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_251
timestamp 1666464484
transform 1 0 24196 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_259
timestamp 1666464484
transform 1 0 24932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_272
timestamp 1666464484
transform 1 0 26128 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1666464484
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_285
timestamp 1666464484
transform 1 0 27324 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1666464484
transform 1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_305
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_311
timestamp 1666464484
transform 1 0 29716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1666464484
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_327
timestamp 1666464484
transform 1 0 31188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_331
timestamp 1666464484
transform 1 0 31556 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1666464484
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_343
timestamp 1666464484
transform 1 0 32660 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_347
timestamp 1666464484
transform 1 0 33028 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_350
timestamp 1666464484
transform 1 0 33304 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_362
timestamp 1666464484
transform 1 0 34408 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_368
timestamp 1666464484
transform 1 0 34960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_375
timestamp 1666464484
transform 1 0 35604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1666464484
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_401
timestamp 1666464484
transform 1 0 37996 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_414
timestamp 1666464484
transform 1 0 39192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_422
timestamp 1666464484
transform 1 0 39928 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_426
timestamp 1666464484
transform 1 0 40296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_430
timestamp 1666464484
transform 1 0 40664 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_436
timestamp 1666464484
transform 1 0 41216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_442
timestamp 1666464484
transform 1 0 41768 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_457
timestamp 1666464484
transform 1 0 43148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_463
timestamp 1666464484
transform 1 0 43700 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_485
timestamp 1666464484
transform 1 0 45724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666464484
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666464484
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_511
timestamp 1666464484
transform 1 0 48116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_526
timestamp 1666464484
transform 1 0 49496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_538
timestamp 1666464484
transform 1 0 50600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_547
timestamp 1666464484
transform 1 0 51428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_551
timestamp 1666464484
transform 1 0 51796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_558
timestamp 1666464484
transform 1 0 52440 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_561
timestamp 1666464484
transform 1 0 52716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_572
timestamp 1666464484
transform 1 0 53728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_580
timestamp 1666464484
transform 1 0 54464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_590
timestamp 1666464484
transform 1 0 55384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_596
timestamp 1666464484
transform 1 0 55936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_602
timestamp 1666464484
transform 1 0 56488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_608
timestamp 1666464484
transform 1 0 57040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_614
timestamp 1666464484
transform 1 0 57592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_617
timestamp 1666464484
transform 1 0 57868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1666464484
transform 1 0 58236 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1666464484
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1666464484
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1666464484
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1666464484
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1666464484
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1666464484
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1666464484
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1666464484
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_259
timestamp 1666464484
transform 1 0 24932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_268
timestamp 1666464484
transform 1 0 25760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1666464484
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_289
timestamp 1666464484
transform 1 0 27692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_300
timestamp 1666464484
transform 1 0 28704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1666464484
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_313
timestamp 1666464484
transform 1 0 29900 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_326
timestamp 1666464484
transform 1 0 31096 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_336
timestamp 1666464484
transform 1 0 32016 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_340
timestamp 1666464484
transform 1 0 32384 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_349
timestamp 1666464484
transform 1 0 33212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1666464484
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_374
timestamp 1666464484
transform 1 0 35512 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_383
timestamp 1666464484
transform 1 0 36340 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_409
timestamp 1666464484
transform 1 0 38732 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_418
timestamp 1666464484
transform 1 0 39560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_429
timestamp 1666464484
transform 1 0 40572 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_439
timestamp 1666464484
transform 1 0 41492 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_456
timestamp 1666464484
transform 1 0 43056 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_460
timestamp 1666464484
transform 1 0 43424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_467
timestamp 1666464484
transform 1 0 44068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_473
timestamp 1666464484
transform 1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_477
timestamp 1666464484
transform 1 0 44988 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_481
timestamp 1666464484
transform 1 0 45356 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_489
timestamp 1666464484
transform 1 0 46092 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_495
timestamp 1666464484
transform 1 0 46644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_507
timestamp 1666464484
transform 1 0 47748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_517
timestamp 1666464484
transform 1 0 48668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_528
timestamp 1666464484
transform 1 0 49680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_533
timestamp 1666464484
transform 1 0 50140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_542
timestamp 1666464484
transform 1 0 50968 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_553
timestamp 1666464484
transform 1 0 51980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_562
timestamp 1666464484
transform 1 0 52808 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_572
timestamp 1666464484
transform 1 0 53728 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_586
timestamp 1666464484
transform 1 0 55016 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_589
timestamp 1666464484
transform 1 0 55292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_596
timestamp 1666464484
transform 1 0 55936 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_602
timestamp 1666464484
transform 1 0 56488 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_608
timestamp 1666464484
transform 1 0 57040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_614
timestamp 1666464484
transform 1 0 57592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_618
timestamp 1666464484
transform 1 0 57960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_622
timestamp 1666464484
transform 1 0 58328 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1666464484
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1666464484
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1666464484
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1666464484
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_255
timestamp 1666464484
transform 1 0 24564 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_260
timestamp 1666464484
transform 1 0 25024 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1666464484
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_291
timestamp 1666464484
transform 1 0 27876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_295
timestamp 1666464484
transform 1 0 28244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_313
timestamp 1666464484
transform 1 0 29900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_324
timestamp 1666464484
transform 1 0 30912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1666464484
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_348
timestamp 1666464484
transform 1 0 33120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_359
timestamp 1666464484
transform 1 0 34132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_365
timestamp 1666464484
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_369
timestamp 1666464484
transform 1 0 35052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_376
timestamp 1666464484
transform 1 0 35696 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1666464484
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_397
timestamp 1666464484
transform 1 0 37628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_408
timestamp 1666464484
transform 1 0 38640 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_418
timestamp 1666464484
transform 1 0 39560 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_427
timestamp 1666464484
transform 1 0 40388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_436
timestamp 1666464484
transform 1 0 41216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_442
timestamp 1666464484
transform 1 0 41768 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_458
timestamp 1666464484
transform 1 0 43240 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_471
timestamp 1666464484
transform 1 0 44436 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_481
timestamp 1666464484
transform 1 0 45356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_487
timestamp 1666464484
transform 1 0 45908 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_496
timestamp 1666464484
transform 1 0 46736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_502
timestamp 1666464484
transform 1 0 47288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_513
timestamp 1666464484
transform 1 0 48300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_517
timestamp 1666464484
transform 1 0 48668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_521
timestamp 1666464484
transform 1 0 49036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_532
timestamp 1666464484
transform 1 0 50048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_538
timestamp 1666464484
transform 1 0 50600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_548
timestamp 1666464484
transform 1 0 51520 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_558
timestamp 1666464484
transform 1 0 52440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_561
timestamp 1666464484
transform 1 0 52716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_570
timestamp 1666464484
transform 1 0 53544 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_586
timestamp 1666464484
transform 1 0 55016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_592
timestamp 1666464484
transform 1 0 55568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_598
timestamp 1666464484
transform 1 0 56120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_604
timestamp 1666464484
transform 1 0 56672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_610
timestamp 1666464484
transform 1 0 57224 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1666464484
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_623
timestamp 1666464484
transform 1 0 58420 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1666464484
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1666464484
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1666464484
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1666464484
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1666464484
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_276
timestamp 1666464484
transform 1 0 26496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_280
timestamp 1666464484
transform 1 0 26864 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_287
timestamp 1666464484
transform 1 0 27508 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_293
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_302
timestamp 1666464484
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_316
timestamp 1666464484
transform 1 0 30176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_322
timestamp 1666464484
transform 1 0 30728 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_326
timestamp 1666464484
transform 1 0 31096 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_340
timestamp 1666464484
transform 1 0 32384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_351
timestamp 1666464484
transform 1 0 33396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_359
timestamp 1666464484
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666464484
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_373
timestamp 1666464484
transform 1 0 35420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_382
timestamp 1666464484
transform 1 0 36248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_386
timestamp 1666464484
transform 1 0 36616 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_390
timestamp 1666464484
transform 1 0 36984 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_405
timestamp 1666464484
transform 1 0 38364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_415
timestamp 1666464484
transform 1 0 39284 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666464484
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_429
timestamp 1666464484
transform 1 0 40572 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_435
timestamp 1666464484
transform 1 0 41124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_441
timestamp 1666464484
transform 1 0 41676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_447
timestamp 1666464484
transform 1 0 42228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_454
timestamp 1666464484
transform 1 0 42872 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_462
timestamp 1666464484
transform 1 0 43608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1666464484
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666464484
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_477
timestamp 1666464484
transform 1 0 44988 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_481
timestamp 1666464484
transform 1 0 45356 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_487
timestamp 1666464484
transform 1 0 45908 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_491
timestamp 1666464484
transform 1 0 46276 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_499
timestamp 1666464484
transform 1 0 47012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_505
timestamp 1666464484
transform 1 0 47564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_514
timestamp 1666464484
transform 1 0 48392 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_522
timestamp 1666464484
transform 1 0 49128 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_530
timestamp 1666464484
transform 1 0 49864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_533
timestamp 1666464484
transform 1 0 50140 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_541
timestamp 1666464484
transform 1 0 50876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_552
timestamp 1666464484
transform 1 0 51888 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_566
timestamp 1666464484
transform 1 0 53176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_575
timestamp 1666464484
transform 1 0 54004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_582
timestamp 1666464484
transform 1 0 54648 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_589
timestamp 1666464484
transform 1 0 55292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_602
timestamp 1666464484
transform 1 0 56488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_608
timestamp 1666464484
transform 1 0 57040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_614
timestamp 1666464484
transform 1 0 57592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_620
timestamp 1666464484
transform 1 0 58144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_624
timestamp 1666464484
transform 1 0 58512 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1666464484
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1666464484
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1666464484
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_245
timestamp 1666464484
transform 1 0 23644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_255
timestamp 1666464484
transform 1 0 24564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_268
timestamp 1666464484
transform 1 0 25760 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1666464484
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_291
timestamp 1666464484
transform 1 0 27876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_299
timestamp 1666464484
transform 1 0 28612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_307
timestamp 1666464484
transform 1 0 29348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_314
timestamp 1666464484
transform 1 0 29992 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_328
timestamp 1666464484
transform 1 0 31280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1666464484
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_346
timestamp 1666464484
transform 1 0 32936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_352
timestamp 1666464484
transform 1 0 33488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_361
timestamp 1666464484
transform 1 0 34316 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_367
timestamp 1666464484
transform 1 0 34868 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_376
timestamp 1666464484
transform 1 0 35696 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1666464484
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_401
timestamp 1666464484
transform 1 0 37996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_405
timestamp 1666464484
transform 1 0 38364 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_412
timestamp 1666464484
transform 1 0 39008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_421
timestamp 1666464484
transform 1 0 39836 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_425
timestamp 1666464484
transform 1 0 40204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_432
timestamp 1666464484
transform 1 0 40848 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1666464484
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_462
timestamp 1666464484
transform 1 0 43608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_475
timestamp 1666464484
transform 1 0 44804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_485
timestamp 1666464484
transform 1 0 45724 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_492
timestamp 1666464484
transform 1 0 46368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_496
timestamp 1666464484
transform 1 0 46736 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_502
timestamp 1666464484
transform 1 0 47288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_514
timestamp 1666464484
transform 1 0 48392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_520
timestamp 1666464484
transform 1 0 48944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_524
timestamp 1666464484
transform 1 0 49312 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_533
timestamp 1666464484
transform 1 0 50140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_544
timestamp 1666464484
transform 1 0 51152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_555
timestamp 1666464484
transform 1 0 52164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1666464484
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_561
timestamp 1666464484
transform 1 0 52716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_572
timestamp 1666464484
transform 1 0 53728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_576
timestamp 1666464484
transform 1 0 54096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_584
timestamp 1666464484
transform 1 0 54832 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_597
timestamp 1666464484
transform 1 0 56028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_603
timestamp 1666464484
transform 1 0 56580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1666464484
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1666464484
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_617
timestamp 1666464484
transform 1 0 57868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_621
timestamp 1666464484
transform 1 0 58236 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1666464484
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1666464484
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1666464484
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1666464484
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_257
timestamp 1666464484
transform 1 0 24748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_263
timestamp 1666464484
transform 1 0 25300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_276
timestamp 1666464484
transform 1 0 26496 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_280
timestamp 1666464484
transform 1 0 26864 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_283
timestamp 1666464484
transform 1 0 27140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_296
timestamp 1666464484
transform 1 0 28336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1666464484
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_314
timestamp 1666464484
transform 1 0 29992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_323
timestamp 1666464484
transform 1 0 30820 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_329
timestamp 1666464484
transform 1 0 31372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_333
timestamp 1666464484
transform 1 0 31740 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_347
timestamp 1666464484
transform 1 0 33028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_356
timestamp 1666464484
transform 1 0 33856 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_362
timestamp 1666464484
transform 1 0 34408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_370
timestamp 1666464484
transform 1 0 35144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_377
timestamp 1666464484
transform 1 0 35788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_383
timestamp 1666464484
transform 1 0 36340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_387
timestamp 1666464484
transform 1 0 36708 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_394
timestamp 1666464484
transform 1 0 37352 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_400
timestamp 1666464484
transform 1 0 37904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_404
timestamp 1666464484
transform 1 0 38272 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_411
timestamp 1666464484
transform 1 0 38916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_417
timestamp 1666464484
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_430
timestamp 1666464484
transform 1 0 40664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_438
timestamp 1666464484
transform 1 0 41400 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_444
timestamp 1666464484
transform 1 0 41952 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_450
timestamp 1666464484
transform 1 0 42504 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_456
timestamp 1666464484
transform 1 0 43056 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_462
timestamp 1666464484
transform 1 0 43608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_466
timestamp 1666464484
transform 1 0 43976 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_473
timestamp 1666464484
transform 1 0 44620 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_477
timestamp 1666464484
transform 1 0 44988 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_492
timestamp 1666464484
transform 1 0 46368 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_500
timestamp 1666464484
transform 1 0 47104 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_507
timestamp 1666464484
transform 1 0 47748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_517
timestamp 1666464484
transform 1 0 48668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_523
timestamp 1666464484
transform 1 0 49220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_529
timestamp 1666464484
transform 1 0 49772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_533
timestamp 1666464484
transform 1 0 50140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_539
timestamp 1666464484
transform 1 0 50692 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_546
timestamp 1666464484
transform 1 0 51336 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_555
timestamp 1666464484
transform 1 0 52164 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_563
timestamp 1666464484
transform 1 0 52900 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_567
timestamp 1666464484
transform 1 0 53268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_579
timestamp 1666464484
transform 1 0 54372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_585
timestamp 1666464484
transform 1 0 54924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_589
timestamp 1666464484
transform 1 0 55292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_593
timestamp 1666464484
transform 1 0 55660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_599
timestamp 1666464484
transform 1 0 56212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_605
timestamp 1666464484
transform 1 0 56764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_611
timestamp 1666464484
transform 1 0 57316 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_617
timestamp 1666464484
transform 1 0 57868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_623
timestamp 1666464484
transform 1 0 58420 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1666464484
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1666464484
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1666464484
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1666464484
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1666464484
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_247
timestamp 1666464484
transform 1 0 23828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_253
timestamp 1666464484
transform 1 0 24380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_263
timestamp 1666464484
transform 1 0 25300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_269
timestamp 1666464484
transform 1 0 25852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_272
timestamp 1666464484
transform 1 0 26128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1666464484
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_290
timestamp 1666464484
transform 1 0 27784 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_296
timestamp 1666464484
transform 1 0 28336 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_304
timestamp 1666464484
transform 1 0 29072 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_316
timestamp 1666464484
transform 1 0 30176 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666464484
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_343
timestamp 1666464484
transform 1 0 32660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_351
timestamp 1666464484
transform 1 0 33396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_360
timestamp 1666464484
transform 1 0 34224 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_366
timestamp 1666464484
transform 1 0 34776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_372
timestamp 1666464484
transform 1 0 35328 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_378
timestamp 1666464484
transform 1 0 35880 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_384
timestamp 1666464484
transform 1 0 36432 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1666464484
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_399
timestamp 1666464484
transform 1 0 37812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_407
timestamp 1666464484
transform 1 0 38548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_413
timestamp 1666464484
transform 1 0 39100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_417
timestamp 1666464484
transform 1 0 39468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_422
timestamp 1666464484
transform 1 0 39928 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_428
timestamp 1666464484
transform 1 0 40480 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_434
timestamp 1666464484
transform 1 0 41032 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_440
timestamp 1666464484
transform 1 0 41584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_446
timestamp 1666464484
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_453
timestamp 1666464484
transform 1 0 42780 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_457
timestamp 1666464484
transform 1 0 43148 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_463
timestamp 1666464484
transform 1 0 43700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_473
timestamp 1666464484
transform 1 0 44620 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_479
timestamp 1666464484
transform 1 0 45172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_483
timestamp 1666464484
transform 1 0 45540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_490
timestamp 1666464484
transform 1 0 46184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_496
timestamp 1666464484
transform 1 0 46736 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_502
timestamp 1666464484
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_513
timestamp 1666464484
transform 1 0 48300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_523
timestamp 1666464484
transform 1 0 49220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_529
timestamp 1666464484
transform 1 0 49772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_535
timestamp 1666464484
transform 1 0 50324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_541
timestamp 1666464484
transform 1 0 50876 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_547
timestamp 1666464484
transform 1 0 51428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_551
timestamp 1666464484
transform 1 0 51796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_558
timestamp 1666464484
transform 1 0 52440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_561
timestamp 1666464484
transform 1 0 52716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_570
timestamp 1666464484
transform 1 0 53544 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_576
timestamp 1666464484
transform 1 0 54096 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_585
timestamp 1666464484
transform 1 0 54924 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_595
timestamp 1666464484
transform 1 0 55844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_602
timestamp 1666464484
transform 1 0 56488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_608
timestamp 1666464484
transform 1 0 57040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_614
timestamp 1666464484
transform 1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_617
timestamp 1666464484
transform 1 0 57868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_621
timestamp 1666464484
transform 1 0 58236 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1666464484
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1666464484
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1666464484
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1666464484
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1666464484
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_259
timestamp 1666464484
transform 1 0 24932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_269
timestamp 1666464484
transform 1 0 25852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_281
timestamp 1666464484
transform 1 0 26956 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_289
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_298
timestamp 1666464484
transform 1 0 28520 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1666464484
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1666464484
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_321
timestamp 1666464484
transform 1 0 30636 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_329
timestamp 1666464484
transform 1 0 31372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_333
timestamp 1666464484
transform 1 0 31740 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_339
timestamp 1666464484
transform 1 0 32292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_343
timestamp 1666464484
transform 1 0 32660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_350
timestamp 1666464484
transform 1 0 33304 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1666464484
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_371
timestamp 1666464484
transform 1 0 35236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_393
timestamp 1666464484
transform 1 0 37260 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_401
timestamp 1666464484
transform 1 0 37996 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_407
timestamp 1666464484
transform 1 0 38548 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1666464484
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_428
timestamp 1666464484
transform 1 0 40480 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_436
timestamp 1666464484
transform 1 0 41216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_441
timestamp 1666464484
transform 1 0 41676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_452
timestamp 1666464484
transform 1 0 42688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_460
timestamp 1666464484
transform 1 0 43424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1666464484
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666464484
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_477
timestamp 1666464484
transform 1 0 44988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_488
timestamp 1666464484
transform 1 0 46000 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_496
timestamp 1666464484
transform 1 0 46736 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_502
timestamp 1666464484
transform 1 0 47288 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_514
timestamp 1666464484
transform 1 0 48392 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_530
timestamp 1666464484
transform 1 0 49864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_533
timestamp 1666464484
transform 1 0 50140 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_537
timestamp 1666464484
transform 1 0 50508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_541
timestamp 1666464484
transform 1 0 50876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_552
timestamp 1666464484
transform 1 0 51888 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_558
timestamp 1666464484
transform 1 0 52440 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_564
timestamp 1666464484
transform 1 0 52992 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_568
timestamp 1666464484
transform 1 0 53360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_575
timestamp 1666464484
transform 1 0 54004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1666464484
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1666464484
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_589
timestamp 1666464484
transform 1 0 55292 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_604
timestamp 1666464484
transform 1 0 56672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_610
timestamp 1666464484
transform 1 0 57224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_616
timestamp 1666464484
transform 1 0 57776 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_622
timestamp 1666464484
transform 1 0 58328 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1666464484
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1666464484
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1666464484
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_252
timestamp 1666464484
transform 1 0 24288 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_260
timestamp 1666464484
transform 1 0 25024 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_266
timestamp 1666464484
transform 1 0 25576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_269
timestamp 1666464484
transform 1 0 25852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1666464484
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_290
timestamp 1666464484
transform 1 0 27784 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_294
timestamp 1666464484
transform 1 0 28152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_304
timestamp 1666464484
transform 1 0 29072 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_318
timestamp 1666464484
transform 1 0 30360 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_324
timestamp 1666464484
transform 1 0 30912 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1666464484
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_346
timestamp 1666464484
transform 1 0 32936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_352
timestamp 1666464484
transform 1 0 33488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_363
timestamp 1666464484
transform 1 0 34500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_376
timestamp 1666464484
transform 1 0 35696 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_382
timestamp 1666464484
transform 1 0 36248 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_390
timestamp 1666464484
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_399
timestamp 1666464484
transform 1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_410
timestamp 1666464484
transform 1 0 38824 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_417
timestamp 1666464484
transform 1 0 39468 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_421
timestamp 1666464484
transform 1 0 39836 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_444
timestamp 1666464484
transform 1 0 41952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_454
timestamp 1666464484
transform 1 0 42872 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_460
timestamp 1666464484
transform 1 0 43424 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_466
timestamp 1666464484
transform 1 0 43976 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_472
timestamp 1666464484
transform 1 0 44528 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_483
timestamp 1666464484
transform 1 0 45540 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_499
timestamp 1666464484
transform 1 0 47012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666464484
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_511
timestamp 1666464484
transform 1 0 48116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_515
timestamp 1666464484
transform 1 0 48484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_520
timestamp 1666464484
transform 1 0 48944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_524
timestamp 1666464484
transform 1 0 49312 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_530
timestamp 1666464484
transform 1 0 49864 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_538
timestamp 1666464484
transform 1 0 50600 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_544
timestamp 1666464484
transform 1 0 51152 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_550
timestamp 1666464484
transform 1 0 51704 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_557
timestamp 1666464484
transform 1 0 52348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_561
timestamp 1666464484
transform 1 0 52716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_566
timestamp 1666464484
transform 1 0 53176 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_574
timestamp 1666464484
transform 1 0 53912 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_582
timestamp 1666464484
transform 1 0 54648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_588
timestamp 1666464484
transform 1 0 55200 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_594
timestamp 1666464484
transform 1 0 55752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_601
timestamp 1666464484
transform 1 0 56396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_607
timestamp 1666464484
transform 1 0 56948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_613
timestamp 1666464484
transform 1 0 57500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_617
timestamp 1666464484
transform 1 0 57868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1666464484
transform 1 0 58236 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1666464484
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1666464484
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_260
timestamp 1666464484
transform 1 0 25024 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_267
timestamp 1666464484
transform 1 0 25668 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_273
timestamp 1666464484
transform 1 0 26220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_276
timestamp 1666464484
transform 1 0 26496 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_282
timestamp 1666464484
transform 1 0 27048 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_291
timestamp 1666464484
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1666464484
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_314
timestamp 1666464484
transform 1 0 29992 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_327
timestamp 1666464484
transform 1 0 31188 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_335
timestamp 1666464484
transform 1 0 31924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_339
timestamp 1666464484
transform 1 0 32292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_347
timestamp 1666464484
transform 1 0 33028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1666464484
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_369
timestamp 1666464484
transform 1 0 35052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_375
timestamp 1666464484
transform 1 0 35604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_381
timestamp 1666464484
transform 1 0 36156 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1666464484
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_399
timestamp 1666464484
transform 1 0 37812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_411
timestamp 1666464484
transform 1 0 38916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_417
timestamp 1666464484
transform 1 0 39468 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_432
timestamp 1666464484
transform 1 0 40848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_438
timestamp 1666464484
transform 1 0 41400 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_444
timestamp 1666464484
transform 1 0 41952 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_450
timestamp 1666464484
transform 1 0 42504 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_457
timestamp 1666464484
transform 1 0 43148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_467
timestamp 1666464484
transform 1 0 44068 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_473
timestamp 1666464484
transform 1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_477
timestamp 1666464484
transform 1 0 44988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_482
timestamp 1666464484
transform 1 0 45448 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_488
timestamp 1666464484
transform 1 0 46000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_494
timestamp 1666464484
transform 1 0 46552 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_500
timestamp 1666464484
transform 1 0 47104 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_508
timestamp 1666464484
transform 1 0 47840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_512
timestamp 1666464484
transform 1 0 48208 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_516
timestamp 1666464484
transform 1 0 48576 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_522
timestamp 1666464484
transform 1 0 49128 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_528
timestamp 1666464484
transform 1 0 49680 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_533
timestamp 1666464484
transform 1 0 50140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_543
timestamp 1666464484
transform 1 0 51060 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_549
timestamp 1666464484
transform 1 0 51612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_558
timestamp 1666464484
transform 1 0 52440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_567
timestamp 1666464484
transform 1 0 53268 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_580
timestamp 1666464484
transform 1 0 54464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_586
timestamp 1666464484
transform 1 0 55016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_589
timestamp 1666464484
transform 1 0 55292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_596
timestamp 1666464484
transform 1 0 55936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_603
timestamp 1666464484
transform 1 0 56580 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_609
timestamp 1666464484
transform 1 0 57132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_615
timestamp 1666464484
transform 1 0 57684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_621
timestamp 1666464484
transform 1 0 58236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1666464484
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1666464484
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1666464484
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1666464484
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1666464484
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1666464484
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1666464484
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_251
timestamp 1666464484
transform 1 0 24196 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1666464484
transform 1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1666464484
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_289
timestamp 1666464484
transform 1 0 27692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_295
timestamp 1666464484
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_299
timestamp 1666464484
transform 1 0 28612 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_307
timestamp 1666464484
transform 1 0 29348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_313
timestamp 1666464484
transform 1 0 29900 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_321
timestamp 1666464484
transform 1 0 30636 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_326
timestamp 1666464484
transform 1 0 31096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1666464484
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_342
timestamp 1666464484
transform 1 0 32568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_348
timestamp 1666464484
transform 1 0 33120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_360
timestamp 1666464484
transform 1 0 34224 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_368
timestamp 1666464484
transform 1 0 34960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_381
timestamp 1666464484
transform 1 0 36156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_388
timestamp 1666464484
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_404
timestamp 1666464484
transform 1 0 38272 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_417
timestamp 1666464484
transform 1 0 39468 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_426
timestamp 1666464484
transform 1 0 40296 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_432
timestamp 1666464484
transform 1 0 40848 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_438
timestamp 1666464484
transform 1 0 41400 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_446
timestamp 1666464484
transform 1 0 42136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_464
timestamp 1666464484
transform 1 0 43792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_468
timestamp 1666464484
transform 1 0 44160 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_477
timestamp 1666464484
transform 1 0 44988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_488
timestamp 1666464484
transform 1 0 46000 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_498
timestamp 1666464484
transform 1 0 46920 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_509
timestamp 1666464484
transform 1 0 47932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_521
timestamp 1666464484
transform 1 0 49036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_530
timestamp 1666464484
transform 1 0 49864 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_546
timestamp 1666464484
transform 1 0 51336 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_558
timestamp 1666464484
transform 1 0 52440 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_561
timestamp 1666464484
transform 1 0 52716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_565
timestamp 1666464484
transform 1 0 53084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_579
timestamp 1666464484
transform 1 0 54372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_588
timestamp 1666464484
transform 1 0 55200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_597
timestamp 1666464484
transform 1 0 56028 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_603
timestamp 1666464484
transform 1 0 56580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1666464484
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1666464484
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_617
timestamp 1666464484
transform 1 0 57868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_621
timestamp 1666464484
transform 1 0 58236 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1666464484
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1666464484
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1666464484
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1666464484
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1666464484
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_257
timestamp 1666464484
transform 1 0 24748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_267
timestamp 1666464484
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_273
timestamp 1666464484
transform 1 0 26220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_279
timestamp 1666464484
transform 1 0 26772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_290
timestamp 1666464484
transform 1 0 27784 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1666464484
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_324
timestamp 1666464484
transform 1 0 30912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_332
timestamp 1666464484
transform 1 0 31648 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_340
timestamp 1666464484
transform 1 0 32384 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_356
timestamp 1666464484
transform 1 0 33856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1666464484
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_371
timestamp 1666464484
transform 1 0 35236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_378
timestamp 1666464484
transform 1 0 35880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_388
timestamp 1666464484
transform 1 0 36800 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_394
timestamp 1666464484
transform 1 0 37352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_404
timestamp 1666464484
transform 1 0 38272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_410
timestamp 1666464484
transform 1 0 38824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1666464484
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_430
timestamp 1666464484
transform 1 0 40664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_436
timestamp 1666464484
transform 1 0 41216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_442
timestamp 1666464484
transform 1 0 41768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_448
timestamp 1666464484
transform 1 0 42320 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_454
timestamp 1666464484
transform 1 0 42872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_463
timestamp 1666464484
transform 1 0 43700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1666464484
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666464484
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_477
timestamp 1666464484
transform 1 0 44988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_483
timestamp 1666464484
transform 1 0 45540 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_491
timestamp 1666464484
transform 1 0 46276 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_500
timestamp 1666464484
transform 1 0 47104 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_506
timestamp 1666464484
transform 1 0 47656 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_520
timestamp 1666464484
transform 1 0 48944 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_524
timestamp 1666464484
transform 1 0 49312 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_528
timestamp 1666464484
transform 1 0 49680 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_533
timestamp 1666464484
transform 1 0 50140 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_544
timestamp 1666464484
transform 1 0 51152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_550
timestamp 1666464484
transform 1 0 51704 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_564
timestamp 1666464484
transform 1 0 52992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_575
timestamp 1666464484
transform 1 0 54004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_585
timestamp 1666464484
transform 1 0 54924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_589
timestamp 1666464484
transform 1 0 55292 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_600
timestamp 1666464484
transform 1 0 56304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_606
timestamp 1666464484
transform 1 0 56856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_612
timestamp 1666464484
transform 1 0 57408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_618
timestamp 1666464484
transform 1 0 57960 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_624
timestamp 1666464484
transform 1 0 58512 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1666464484
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1666464484
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1666464484
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1666464484
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1666464484
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1666464484
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_245
timestamp 1666464484
transform 1 0 23644 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_248
timestamp 1666464484
transform 1 0 23920 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_255
timestamp 1666464484
transform 1 0 24564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_265
timestamp 1666464484
transform 1 0 25484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1666464484
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_293
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_299
timestamp 1666464484
transform 1 0 28612 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_306
timestamp 1666464484
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_313
timestamp 1666464484
transform 1 0 29900 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_321
timestamp 1666464484
transform 1 0 30636 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1666464484
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666464484
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_346
timestamp 1666464484
transform 1 0 32936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_356
timestamp 1666464484
transform 1 0 33856 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_362
timestamp 1666464484
transform 1 0 34408 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_377
timestamp 1666464484
transform 1 0 35788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1666464484
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666464484
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_397
timestamp 1666464484
transform 1 0 37628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_404
timestamp 1666464484
transform 1 0 38272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_408
timestamp 1666464484
transform 1 0 38640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_415
timestamp 1666464484
transform 1 0 39284 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_429
timestamp 1666464484
transform 1 0 40572 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_435
timestamp 1666464484
transform 1 0 41124 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_441
timestamp 1666464484
transform 1 0 41676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1666464484
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_458
timestamp 1666464484
transform 1 0 43240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_465
timestamp 1666464484
transform 1 0 43884 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_475
timestamp 1666464484
transform 1 0 44804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_481
timestamp 1666464484
transform 1 0 45356 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_492
timestamp 1666464484
transform 1 0 46368 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_500
timestamp 1666464484
transform 1 0 47104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_511
timestamp 1666464484
transform 1 0 48116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_519
timestamp 1666464484
transform 1 0 48852 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_528
timestamp 1666464484
transform 1 0 49680 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_541
timestamp 1666464484
transform 1 0 50876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_547
timestamp 1666464484
transform 1 0 51428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_558
timestamp 1666464484
transform 1 0 52440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_561
timestamp 1666464484
transform 1 0 52716 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_569
timestamp 1666464484
transform 1 0 53452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_575
timestamp 1666464484
transform 1 0 54004 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_581
timestamp 1666464484
transform 1 0 54556 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_587
timestamp 1666464484
transform 1 0 55108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_595
timestamp 1666464484
transform 1 0 55844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_601
timestamp 1666464484
transform 1 0 56396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_607
timestamp 1666464484
transform 1 0 56948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_613
timestamp 1666464484
transform 1 0 57500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_617
timestamp 1666464484
transform 1 0 57868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_621
timestamp 1666464484
transform 1 0 58236 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1666464484
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1666464484
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1666464484
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1666464484
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_245
timestamp 1666464484
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1666464484
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_263
timestamp 1666464484
transform 1 0 25300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_273
timestamp 1666464484
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_282
timestamp 1666464484
transform 1 0 27048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_293
timestamp 1666464484
transform 1 0 28060 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1666464484
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_316
timestamp 1666464484
transform 1 0 30176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_320
timestamp 1666464484
transform 1 0 30544 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_329
timestamp 1666464484
transform 1 0 31372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_335
timestamp 1666464484
transform 1 0 31924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_341
timestamp 1666464484
transform 1 0 32476 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_347
timestamp 1666464484
transform 1 0 33028 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_350
timestamp 1666464484
transform 1 0 33304 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1666464484
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_369
timestamp 1666464484
transform 1 0 35052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_375
timestamp 1666464484
transform 1 0 35604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_381
timestamp 1666464484
transform 1 0 36156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_387
timestamp 1666464484
transform 1 0 36708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_397
timestamp 1666464484
transform 1 0 37628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_404
timestamp 1666464484
transform 1 0 38272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_410
timestamp 1666464484
transform 1 0 38824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1666464484
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_432
timestamp 1666464484
transform 1 0 40848 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_438
timestamp 1666464484
transform 1 0 41400 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_451
timestamp 1666464484
transform 1 0 42596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_458
timestamp 1666464484
transform 1 0 43240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_470
timestamp 1666464484
transform 1 0 44344 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_477
timestamp 1666464484
transform 1 0 44988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_481
timestamp 1666464484
transform 1 0 45356 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_493
timestamp 1666464484
transform 1 0 46460 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_501
timestamp 1666464484
transform 1 0 47196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_509
timestamp 1666464484
transform 1 0 47932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_518
timestamp 1666464484
transform 1 0 48760 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_528
timestamp 1666464484
transform 1 0 49680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_533
timestamp 1666464484
transform 1 0 50140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_541
timestamp 1666464484
transform 1 0 50876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_551
timestamp 1666464484
transform 1 0 51796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_557
timestamp 1666464484
transform 1 0 52348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_563
timestamp 1666464484
transform 1 0 52900 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_569
timestamp 1666464484
transform 1 0 53452 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_573
timestamp 1666464484
transform 1 0 53820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_583
timestamp 1666464484
transform 1 0 54740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1666464484
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_589
timestamp 1666464484
transform 1 0 55292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_599
timestamp 1666464484
transform 1 0 56212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_605
timestamp 1666464484
transform 1 0 56764 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_611
timestamp 1666464484
transform 1 0 57316 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_623
timestamp 1666464484
transform 1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1666464484
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1666464484
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1666464484
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1666464484
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_252
timestamp 1666464484
transform 1 0 24288 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_260
timestamp 1666464484
transform 1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_269
timestamp 1666464484
transform 1 0 25852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1666464484
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_287
timestamp 1666464484
transform 1 0 27508 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_295
timestamp 1666464484
transform 1 0 28244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_302
timestamp 1666464484
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_306
timestamp 1666464484
transform 1 0 29256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_314
timestamp 1666464484
transform 1 0 29992 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_326
timestamp 1666464484
transform 1 0 31096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1666464484
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_345
timestamp 1666464484
transform 1 0 32844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_355
timestamp 1666464484
transform 1 0 33764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_361
timestamp 1666464484
transform 1 0 34316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_368
timestamp 1666464484
transform 1 0 34960 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_374
timestamp 1666464484
transform 1 0 35512 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_382
timestamp 1666464484
transform 1 0 36248 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_386
timestamp 1666464484
transform 1 0 36616 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1666464484
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_400
timestamp 1666464484
transform 1 0 37904 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_406
timestamp 1666464484
transform 1 0 38456 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_415
timestamp 1666464484
transform 1 0 39284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_424
timestamp 1666464484
transform 1 0 40112 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_434
timestamp 1666464484
transform 1 0 41032 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_442
timestamp 1666464484
transform 1 0 41768 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_453
timestamp 1666464484
transform 1 0 42780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_457
timestamp 1666464484
transform 1 0 43148 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_463
timestamp 1666464484
transform 1 0 43700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_471
timestamp 1666464484
transform 1 0 44436 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_475
timestamp 1666464484
transform 1 0 44804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_484
timestamp 1666464484
transform 1 0 45632 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_492
timestamp 1666464484
transform 1 0 46368 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_502
timestamp 1666464484
transform 1 0 47288 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_509
timestamp 1666464484
transform 1 0 47932 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_517
timestamp 1666464484
transform 1 0 48668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_523
timestamp 1666464484
transform 1 0 49220 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_531
timestamp 1666464484
transform 1 0 49956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_539
timestamp 1666464484
transform 1 0 50692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_546
timestamp 1666464484
transform 1 0 51336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_554
timestamp 1666464484
transform 1 0 52072 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_558
timestamp 1666464484
transform 1 0 52440 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_561
timestamp 1666464484
transform 1 0 52716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_571
timestamp 1666464484
transform 1 0 53636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_582
timestamp 1666464484
transform 1 0 54648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_588
timestamp 1666464484
transform 1 0 55200 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1666464484
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1666464484
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_617
timestamp 1666464484
transform 1 0 57868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_621
timestamp 1666464484
transform 1 0 58236 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1666464484
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1666464484
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1666464484
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1666464484
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_229
timestamp 1666464484
transform 1 0 22172 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1666464484
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1666464484
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_264
timestamp 1666464484
transform 1 0 25392 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_268
timestamp 1666464484
transform 1 0 25760 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1666464484
transform 1 0 26036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1666464484
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1666464484
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_297
timestamp 1666464484
transform 1 0 28428 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_303
timestamp 1666464484
transform 1 0 28980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666464484
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_321
timestamp 1666464484
transform 1 0 30636 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_335
timestamp 1666464484
transform 1 0 31924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_347
timestamp 1666464484
transform 1 0 33028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1666464484
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_375
timestamp 1666464484
transform 1 0 35604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_381
timestamp 1666464484
transform 1 0 36156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_390
timestamp 1666464484
transform 1 0 36984 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_394
timestamp 1666464484
transform 1 0 37352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_401
timestamp 1666464484
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666464484
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666464484
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_431
timestamp 1666464484
transform 1 0 40756 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_437
timestamp 1666464484
transform 1 0 41308 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_444
timestamp 1666464484
transform 1 0 41952 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_454
timestamp 1666464484
transform 1 0 42872 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_460
timestamp 1666464484
transform 1 0 43424 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_466
timestamp 1666464484
transform 1 0 43976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_472
timestamp 1666464484
transform 1 0 44528 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_477
timestamp 1666464484
transform 1 0 44988 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_483
timestamp 1666464484
transform 1 0 45540 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_492
timestamp 1666464484
transform 1 0 46368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_496
timestamp 1666464484
transform 1 0 46736 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_505
timestamp 1666464484
transform 1 0 47564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_509
timestamp 1666464484
transform 1 0 47932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_516
timestamp 1666464484
transform 1 0 48576 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_524
timestamp 1666464484
transform 1 0 49312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_530
timestamp 1666464484
transform 1 0 49864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_533
timestamp 1666464484
transform 1 0 50140 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_539
timestamp 1666464484
transform 1 0 50692 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_548
timestamp 1666464484
transform 1 0 51520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_560
timestamp 1666464484
transform 1 0 52624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_571
timestamp 1666464484
transform 1 0 53636 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_580
timestamp 1666464484
transform 1 0 54464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_586
timestamp 1666464484
transform 1 0 55016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_589
timestamp 1666464484
transform 1 0 55292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_594
timestamp 1666464484
transform 1 0 55752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_600
timestamp 1666464484
transform 1 0 56304 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_606
timestamp 1666464484
transform 1 0 56856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_612
timestamp 1666464484
transform 1 0 57408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_618
timestamp 1666464484
transform 1 0 57960 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_624
timestamp 1666464484
transform 1 0 58512 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1666464484
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1666464484
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1666464484
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1666464484
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1666464484
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_237
timestamp 1666464484
transform 1 0 22908 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_254
timestamp 1666464484
transform 1 0 24472 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_260
timestamp 1666464484
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_269
timestamp 1666464484
transform 1 0 25852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1666464484
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_290
timestamp 1666464484
transform 1 0 27784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1666464484
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_306
timestamp 1666464484
transform 1 0 29256 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_319
timestamp 1666464484
transform 1 0 30452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1666464484
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_341
timestamp 1666464484
transform 1 0 32476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_347
timestamp 1666464484
transform 1 0 33028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_353
timestamp 1666464484
transform 1 0 33580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_359
timestamp 1666464484
transform 1 0 34132 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_368
timestamp 1666464484
transform 1 0 34960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_375
timestamp 1666464484
transform 1 0 35604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_386
timestamp 1666464484
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_400
timestamp 1666464484
transform 1 0 37904 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_406
timestamp 1666464484
transform 1 0 38456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_410
timestamp 1666464484
transform 1 0 38824 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_418
timestamp 1666464484
transform 1 0 39560 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_424
timestamp 1666464484
transform 1 0 40112 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_428
timestamp 1666464484
transform 1 0 40480 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_442
timestamp 1666464484
transform 1 0 41768 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_455
timestamp 1666464484
transform 1 0 42964 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_466
timestamp 1666464484
transform 1 0 43976 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_472
timestamp 1666464484
transform 1 0 44528 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_480
timestamp 1666464484
transform 1 0 45264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_491
timestamp 1666464484
transform 1 0 46276 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_495
timestamp 1666464484
transform 1 0 46644 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_501
timestamp 1666464484
transform 1 0 47196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_512
timestamp 1666464484
transform 1 0 48208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_524
timestamp 1666464484
transform 1 0 49312 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_536
timestamp 1666464484
transform 1 0 50416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_545
timestamp 1666464484
transform 1 0 51244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_558
timestamp 1666464484
transform 1 0 52440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_561
timestamp 1666464484
transform 1 0 52716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_568
timestamp 1666464484
transform 1 0 53360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_572
timestamp 1666464484
transform 1 0 53728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_580
timestamp 1666464484
transform 1 0 54464 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_610
timestamp 1666464484
transform 1 0 57224 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_617
timestamp 1666464484
transform 1 0 57868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_621
timestamp 1666464484
transform 1 0 58236 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1666464484
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1666464484
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1666464484
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1666464484
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1666464484
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_235
timestamp 1666464484
transform 1 0 22724 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_241
timestamp 1666464484
transform 1 0 23276 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1666464484
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666464484
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_259
timestamp 1666464484
transform 1 0 24932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_263
timestamp 1666464484
transform 1 0 25300 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_266
timestamp 1666464484
transform 1 0 25576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_270
timestamp 1666464484
transform 1 0 25944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_278
timestamp 1666464484
transform 1 0 26680 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_286
timestamp 1666464484
transform 1 0 27416 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_293
timestamp 1666464484
transform 1 0 28060 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1666464484
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_318
timestamp 1666464484
transform 1 0 30360 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_324
timestamp 1666464484
transform 1 0 30912 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_329
timestamp 1666464484
transform 1 0 31372 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_342
timestamp 1666464484
transform 1 0 32568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_350
timestamp 1666464484
transform 1 0 33304 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_358
timestamp 1666464484
transform 1 0 34040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1666464484
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_376
timestamp 1666464484
transform 1 0 35696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_387
timestamp 1666464484
transform 1 0 36708 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1666464484
transform 1 0 37260 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_401
timestamp 1666464484
transform 1 0 37996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_405
timestamp 1666464484
transform 1 0 38364 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_415
timestamp 1666464484
transform 1 0 39284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1666464484
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_425
timestamp 1666464484
transform 1 0 40204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_437
timestamp 1666464484
transform 1 0 41308 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_445
timestamp 1666464484
transform 1 0 42044 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_451
timestamp 1666464484
transform 1 0 42596 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_461
timestamp 1666464484
transform 1 0 43516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_471
timestamp 1666464484
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666464484
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_477
timestamp 1666464484
transform 1 0 44988 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_484
timestamp 1666464484
transform 1 0 45632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_488
timestamp 1666464484
transform 1 0 46000 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_496
timestamp 1666464484
transform 1 0 46736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_509
timestamp 1666464484
transform 1 0 47932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_515
timestamp 1666464484
transform 1 0 48484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_521
timestamp 1666464484
transform 1 0 49036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_530
timestamp 1666464484
transform 1 0 49864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_533
timestamp 1666464484
transform 1 0 50140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_541
timestamp 1666464484
transform 1 0 50876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_547
timestamp 1666464484
transform 1 0 51428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_551
timestamp 1666464484
transform 1 0 51796 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_558
timestamp 1666464484
transform 1 0 52440 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_568
timestamp 1666464484
transform 1 0 53360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_574
timestamp 1666464484
transform 1 0 53912 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_580
timestamp 1666464484
transform 1 0 54464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_586
timestamp 1666464484
transform 1 0 55016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_589
timestamp 1666464484
transform 1 0 55292 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_597
timestamp 1666464484
transform 1 0 56028 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_603
timestamp 1666464484
transform 1 0 56580 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_609
timestamp 1666464484
transform 1 0 57132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_615
timestamp 1666464484
transform 1 0 57684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_621
timestamp 1666464484
transform 1 0 58236 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1666464484
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1666464484
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1666464484
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1666464484
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_247
timestamp 1666464484
transform 1 0 23828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_260
timestamp 1666464484
transform 1 0 25024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_266
timestamp 1666464484
transform 1 0 25576 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_270
timestamp 1666464484
transform 1 0 25944 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1666464484
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_289
timestamp 1666464484
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1666464484
transform 1 0 28244 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_301
timestamp 1666464484
transform 1 0 28796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_307
timestamp 1666464484
transform 1 0 29348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_317
timestamp 1666464484
transform 1 0 30268 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1666464484
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_350
timestamp 1666464484
transform 1 0 33304 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_358
timestamp 1666464484
transform 1 0 34040 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_370
timestamp 1666464484
transform 1 0 35144 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_381
timestamp 1666464484
transform 1 0 36156 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1666464484
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_404
timestamp 1666464484
transform 1 0 38272 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_410
timestamp 1666464484
transform 1 0 38824 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_422
timestamp 1666464484
transform 1 0 39928 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_431
timestamp 1666464484
transform 1 0 40756 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_443
timestamp 1666464484
transform 1 0 41860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1666464484
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_456
timestamp 1666464484
transform 1 0 43056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_460
timestamp 1666464484
transform 1 0 43424 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_464
timestamp 1666464484
transform 1 0 43792 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_475
timestamp 1666464484
transform 1 0 44804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_492
timestamp 1666464484
transform 1 0 46368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_499
timestamp 1666464484
transform 1 0 47012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666464484
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_510
timestamp 1666464484
transform 1 0 48024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_514
timestamp 1666464484
transform 1 0 48392 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_522
timestamp 1666464484
transform 1 0 49128 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_528
timestamp 1666464484
transform 1 0 49680 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_532
timestamp 1666464484
transform 1 0 50048 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_551
timestamp 1666464484
transform 1 0 51796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_557
timestamp 1666464484
transform 1 0 52348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_561
timestamp 1666464484
transform 1 0 52716 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_565
timestamp 1666464484
transform 1 0 53084 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_578
timestamp 1666464484
transform 1 0 54280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_582
timestamp 1666464484
transform 1 0 54648 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_589
timestamp 1666464484
transform 1 0 55292 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_595
timestamp 1666464484
transform 1 0 55844 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_599
timestamp 1666464484
transform 1 0 56212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_605
timestamp 1666464484
transform 1 0 56764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_611
timestamp 1666464484
transform 1 0 57316 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1666464484
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_617
timestamp 1666464484
transform 1 0 57868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1666464484
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1666464484
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1666464484
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1666464484
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_229
timestamp 1666464484
transform 1 0 22172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1666464484
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_257
timestamp 1666464484
transform 1 0 24748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_269
timestamp 1666464484
transform 1 0 25852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_292
timestamp 1666464484
transform 1 0 27968 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_300
timestamp 1666464484
transform 1 0 28704 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1666464484
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_319
timestamp 1666464484
transform 1 0 30452 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_325
timestamp 1666464484
transform 1 0 31004 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_329
timestamp 1666464484
transform 1 0 31372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_336
timestamp 1666464484
transform 1 0 32016 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_353
timestamp 1666464484
transform 1 0 33580 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1666464484
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_377
timestamp 1666464484
transform 1 0 35788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_385
timestamp 1666464484
transform 1 0 36524 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_395
timestamp 1666464484
transform 1 0 37444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_408
timestamp 1666464484
transform 1 0 38640 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_412
timestamp 1666464484
transform 1 0 39008 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1666464484
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_429
timestamp 1666464484
transform 1 0 40572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_459
timestamp 1666464484
transform 1 0 43332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1666464484
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666464484
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_477
timestamp 1666464484
transform 1 0 44988 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_498
timestamp 1666464484
transform 1 0 46920 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_516
timestamp 1666464484
transform 1 0 48576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1666464484
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_533
timestamp 1666464484
transform 1 0 50140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_540
timestamp 1666464484
transform 1 0 50784 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_551
timestamp 1666464484
transform 1 0 51796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_563
timestamp 1666464484
transform 1 0 52900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_573
timestamp 1666464484
transform 1 0 53820 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_579
timestamp 1666464484
transform 1 0 54372 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_584
timestamp 1666464484
transform 1 0 54832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_589
timestamp 1666464484
transform 1 0 55292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_598
timestamp 1666464484
transform 1 0 56120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_606
timestamp 1666464484
transform 1 0 56856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_612
timestamp 1666464484
transform 1 0 57408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_618
timestamp 1666464484
transform 1 0 57960 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_624
timestamp 1666464484
transform 1 0 58512 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1666464484
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1666464484
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1666464484
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1666464484
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_234
timestamp 1666464484
transform 1 0 22632 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_246
timestamp 1666464484
transform 1 0 23736 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_249
timestamp 1666464484
transform 1 0 24012 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_260
timestamp 1666464484
transform 1 0 25024 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_268
timestamp 1666464484
transform 1 0 25760 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1666464484
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_287
timestamp 1666464484
transform 1 0 27508 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1666464484
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_301
timestamp 1666464484
transform 1 0 28796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_309
timestamp 1666464484
transform 1 0 29532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_315
timestamp 1666464484
transform 1 0 30084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_319
timestamp 1666464484
transform 1 0 30452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_328
timestamp 1666464484
transform 1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_344
timestamp 1666464484
transform 1 0 32752 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_352
timestamp 1666464484
transform 1 0 33488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_359
timestamp 1666464484
transform 1 0 34132 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_372
timestamp 1666464484
transform 1 0 35328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1666464484
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666464484
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_399
timestamp 1666464484
transform 1 0 37812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_407
timestamp 1666464484
transform 1 0 38548 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_413
timestamp 1666464484
transform 1 0 39100 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_421
timestamp 1666464484
transform 1 0 39836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_426
timestamp 1666464484
transform 1 0 40296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_436
timestamp 1666464484
transform 1 0 41216 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1666464484
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_456
timestamp 1666464484
transform 1 0 43056 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_465
timestamp 1666464484
transform 1 0 43884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_476
timestamp 1666464484
transform 1 0 44896 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_482
timestamp 1666464484
transform 1 0 45448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_486
timestamp 1666464484
transform 1 0 45816 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_490
timestamp 1666464484
transform 1 0 46184 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_502
timestamp 1666464484
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_509
timestamp 1666464484
transform 1 0 47932 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_515
timestamp 1666464484
transform 1 0 48484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_537
timestamp 1666464484
transform 1 0 50508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_549
timestamp 1666464484
transform 1 0 51612 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_557
timestamp 1666464484
transform 1 0 52348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_561
timestamp 1666464484
transform 1 0 52716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_569
timestamp 1666464484
transform 1 0 53452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_576
timestamp 1666464484
transform 1 0 54096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_585
timestamp 1666464484
transform 1 0 54924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_591
timestamp 1666464484
transform 1 0 55476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_602
timestamp 1666464484
transform 1 0 56488 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_608
timestamp 1666464484
transform 1 0 57040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_614
timestamp 1666464484
transform 1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_617
timestamp 1666464484
transform 1 0 57868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1666464484
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1666464484
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1666464484
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1666464484
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1666464484
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_233
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_239
timestamp 1666464484
transform 1 0 23092 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_242
timestamp 1666464484
transform 1 0 23368 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1666464484
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_262
timestamp 1666464484
transform 1 0 25208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_268
timestamp 1666464484
transform 1 0 25760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_277
timestamp 1666464484
transform 1 0 26588 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_283
timestamp 1666464484
transform 1 0 27140 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_288
timestamp 1666464484
transform 1 0 27600 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_297
timestamp 1666464484
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1666464484
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_321
timestamp 1666464484
transform 1 0 30636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_329
timestamp 1666464484
transform 1 0 31372 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_337
timestamp 1666464484
transform 1 0 32108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_349
timestamp 1666464484
transform 1 0 33212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1666464484
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666464484
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_372
timestamp 1666464484
transform 1 0 35328 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_384
timestamp 1666464484
transform 1 0 36432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_396
timestamp 1666464484
transform 1 0 37536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_403
timestamp 1666464484
transform 1 0 38180 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_409
timestamp 1666464484
transform 1 0 38732 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_415
timestamp 1666464484
transform 1 0 39284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666464484
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_427
timestamp 1666464484
transform 1 0 40388 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_430
timestamp 1666464484
transform 1 0 40664 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_442
timestamp 1666464484
transform 1 0 41768 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_450
timestamp 1666464484
transform 1 0 42504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_454
timestamp 1666464484
transform 1 0 42872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_466
timestamp 1666464484
transform 1 0 43976 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1666464484
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_477
timestamp 1666464484
transform 1 0 44988 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_486
timestamp 1666464484
transform 1 0 45816 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_500
timestamp 1666464484
transform 1 0 47104 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_506
timestamp 1666464484
transform 1 0 47656 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_517
timestamp 1666464484
transform 1 0 48668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_525
timestamp 1666464484
transform 1 0 49404 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_530
timestamp 1666464484
transform 1 0 49864 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_533
timestamp 1666464484
transform 1 0 50140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_543
timestamp 1666464484
transform 1 0 51060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_559
timestamp 1666464484
transform 1 0 52532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_563
timestamp 1666464484
transform 1 0 52900 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_569
timestamp 1666464484
transform 1 0 53452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_578
timestamp 1666464484
transform 1 0 54280 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_584
timestamp 1666464484
transform 1 0 54832 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_589
timestamp 1666464484
transform 1 0 55292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_600
timestamp 1666464484
transform 1 0 56304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_606
timestamp 1666464484
transform 1 0 56856 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_612
timestamp 1666464484
transform 1 0 57408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_618
timestamp 1666464484
transform 1 0 57960 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_624
timestamp 1666464484
transform 1 0 58512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_9
timestamp 1666464484
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1666464484
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1666464484
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1666464484
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1666464484
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1666464484
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1666464484
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_250
timestamp 1666464484
transform 1 0 24104 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_261
timestamp 1666464484
transform 1 0 25116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_269
timestamp 1666464484
transform 1 0 25852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1666464484
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1666464484
transform 1 0 27416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_297
timestamp 1666464484
transform 1 0 28428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_305
timestamp 1666464484
transform 1 0 29164 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_315
timestamp 1666464484
transform 1 0 30084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_322
timestamp 1666464484
transform 1 0 30728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1666464484
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1666464484
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1666464484
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_373
timestamp 1666464484
transform 1 0 35420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_383
timestamp 1666464484
transform 1 0 36340 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_387
timestamp 1666464484
transform 1 0 36708 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1666464484
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_399
timestamp 1666464484
transform 1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_406
timestamp 1666464484
transform 1 0 38456 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_414
timestamp 1666464484
transform 1 0 39192 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_421
timestamp 1666464484
transform 1 0 39836 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_433
timestamp 1666464484
transform 1 0 40940 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_439
timestamp 1666464484
transform 1 0 41492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1666464484
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_454
timestamp 1666464484
transform 1 0 42872 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_460
timestamp 1666464484
transform 1 0 43424 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_468
timestamp 1666464484
transform 1 0 44160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_479
timestamp 1666464484
transform 1 0 45172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_483
timestamp 1666464484
transform 1 0 45540 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_493
timestamp 1666464484
transform 1 0 46460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_499
timestamp 1666464484
transform 1 0 47012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666464484
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_509
timestamp 1666464484
transform 1 0 47932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_516
timestamp 1666464484
transform 1 0 48576 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_523
timestamp 1666464484
transform 1 0 49220 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_536
timestamp 1666464484
transform 1 0 50416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_542
timestamp 1666464484
transform 1 0 50968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_548
timestamp 1666464484
transform 1 0 51520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_554
timestamp 1666464484
transform 1 0 52072 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_561
timestamp 1666464484
transform 1 0 52716 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_567
timestamp 1666464484
transform 1 0 53268 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_575
timestamp 1666464484
transform 1 0 54004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_581
timestamp 1666464484
transform 1 0 54556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_585
timestamp 1666464484
transform 1 0 54924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_589
timestamp 1666464484
transform 1 0 55292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_598
timestamp 1666464484
transform 1 0 56120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_604
timestamp 1666464484
transform 1 0 56672 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_610
timestamp 1666464484
transform 1 0 57224 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_617
timestamp 1666464484
transform 1 0 57868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_621
timestamp 1666464484
transform 1 0 58236 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1666464484
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1666464484
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1666464484
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1666464484
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_223
timestamp 1666464484
transform 1 0 21620 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_230
timestamp 1666464484
transform 1 0 22264 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_238
timestamp 1666464484
transform 1 0 23000 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1666464484
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_257
timestamp 1666464484
transform 1 0 24748 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_263
timestamp 1666464484
transform 1 0 25300 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_269
timestamp 1666464484
transform 1 0 25852 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_278
timestamp 1666464484
transform 1 0 26680 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_290
timestamp 1666464484
transform 1 0 27784 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_302
timestamp 1666464484
transform 1 0 28888 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1666464484
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_315
timestamp 1666464484
transform 1 0 30084 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_323
timestamp 1666464484
transform 1 0 30820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_337
timestamp 1666464484
transform 1 0 32108 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_348
timestamp 1666464484
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1666464484
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_373
timestamp 1666464484
transform 1 0 35420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_382
timestamp 1666464484
transform 1 0 36248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_391
timestamp 1666464484
transform 1 0 37076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_404
timestamp 1666464484
transform 1 0 38272 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 1666464484
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_432
timestamp 1666464484
transform 1 0 40848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_443
timestamp 1666464484
transform 1 0 41860 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_451
timestamp 1666464484
transform 1 0 42596 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_462
timestamp 1666464484
transform 1 0 43608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_466
timestamp 1666464484
transform 1 0 43976 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1666464484
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1666464484
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_477
timestamp 1666464484
transform 1 0 44988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_481
timestamp 1666464484
transform 1 0 45356 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_489
timestamp 1666464484
transform 1 0 46092 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_499
timestamp 1666464484
transform 1 0 47012 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_506
timestamp 1666464484
transform 1 0 47656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1666464484
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_518
timestamp 1666464484
transform 1 0 48760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_524
timestamp 1666464484
transform 1 0 49312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_530
timestamp 1666464484
transform 1 0 49864 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_533
timestamp 1666464484
transform 1 0 50140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_544
timestamp 1666464484
transform 1 0 51152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_548
timestamp 1666464484
transform 1 0 51520 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_562
timestamp 1666464484
transform 1 0 52808 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_583
timestamp 1666464484
transform 1 0 54740 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1666464484
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_589
timestamp 1666464484
transform 1 0 55292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_599
timestamp 1666464484
transform 1 0 56212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_605
timestamp 1666464484
transform 1 0 56764 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_611
timestamp 1666464484
transform 1 0 57316 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_623
timestamp 1666464484
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1666464484
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1666464484
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_247
timestamp 1666464484
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_260
timestamp 1666464484
transform 1 0 25024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_267
timestamp 1666464484
transform 1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1666464484
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_285
timestamp 1666464484
transform 1 0 27324 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_296
timestamp 1666464484
transform 1 0 28336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_303
timestamp 1666464484
transform 1 0 28980 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_316
timestamp 1666464484
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_328
timestamp 1666464484
transform 1 0 31280 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1666464484
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_347
timestamp 1666464484
transform 1 0 33028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_356
timestamp 1666464484
transform 1 0 33856 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_368
timestamp 1666464484
transform 1 0 34960 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_380
timestamp 1666464484
transform 1 0 36064 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1666464484
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_402
timestamp 1666464484
transform 1 0 38088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_414
timestamp 1666464484
transform 1 0 39192 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_417
timestamp 1666464484
transform 1 0 39468 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_426
timestamp 1666464484
transform 1 0 40296 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_434
timestamp 1666464484
transform 1 0 41032 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_438
timestamp 1666464484
transform 1 0 41400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1666464484
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_454
timestamp 1666464484
transform 1 0 42872 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_467
timestamp 1666464484
transform 1 0 44068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_473
timestamp 1666464484
transform 1 0 44620 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_479
timestamp 1666464484
transform 1 0 45172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_483
timestamp 1666464484
transform 1 0 45540 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_491
timestamp 1666464484
transform 1 0 46276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1666464484
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666464484
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_509
timestamp 1666464484
transform 1 0 47932 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_513
timestamp 1666464484
transform 1 0 48300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_525
timestamp 1666464484
transform 1 0 49404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_539
timestamp 1666464484
transform 1 0 50692 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_545
timestamp 1666464484
transform 1 0 51244 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_555
timestamp 1666464484
transform 1 0 52164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1666464484
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_561
timestamp 1666464484
transform 1 0 52716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_569
timestamp 1666464484
transform 1 0 53452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_575
timestamp 1666464484
transform 1 0 54004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_581
timestamp 1666464484
transform 1 0 54556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_585
timestamp 1666464484
transform 1 0 54924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_595
timestamp 1666464484
transform 1 0 55844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_610
timestamp 1666464484
transform 1 0 57224 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_617
timestamp 1666464484
transform 1 0 57868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_621
timestamp 1666464484
transform 1 0 58236 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1666464484
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1666464484
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1666464484
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_233
timestamp 1666464484
transform 1 0 22540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_241
timestamp 1666464484
transform 1 0 23276 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1666464484
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_268
timestamp 1666464484
transform 1 0 25760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_283
timestamp 1666464484
transform 1 0 27140 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_291
timestamp 1666464484
transform 1 0 27876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_300
timestamp 1666464484
transform 1 0 28704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1666464484
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_316
timestamp 1666464484
transform 1 0 30176 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_328
timestamp 1666464484
transform 1 0 31280 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1666464484
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_345
timestamp 1666464484
transform 1 0 32844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_349
timestamp 1666464484
transform 1 0 33212 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_354
timestamp 1666464484
transform 1 0 33672 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1666464484
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_376
timestamp 1666464484
transform 1 0 35696 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_393
timestamp 1666464484
transform 1 0 37260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_404
timestamp 1666464484
transform 1 0 38272 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_408
timestamp 1666464484
transform 1 0 38640 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_415
timestamp 1666464484
transform 1 0 39284 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666464484
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_428
timestamp 1666464484
transform 1 0 40480 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_434
timestamp 1666464484
transform 1 0 41032 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_448
timestamp 1666464484
transform 1 0 42320 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_452
timestamp 1666464484
transform 1 0 42688 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_465
timestamp 1666464484
transform 1 0 43884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1666464484
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_477
timestamp 1666464484
transform 1 0 44988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_488
timestamp 1666464484
transform 1 0 46000 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_492
timestamp 1666464484
transform 1 0 46368 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_499
timestamp 1666464484
transform 1 0 47012 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_510
timestamp 1666464484
transform 1 0 48024 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_524
timestamp 1666464484
transform 1 0 49312 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_533
timestamp 1666464484
transform 1 0 50140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_545
timestamp 1666464484
transform 1 0 51244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_558
timestamp 1666464484
transform 1 0 52440 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_572
timestamp 1666464484
transform 1 0 53728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_582
timestamp 1666464484
transform 1 0 54648 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_589
timestamp 1666464484
transform 1 0 55292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_595
timestamp 1666464484
transform 1 0 55844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_605
timestamp 1666464484
transform 1 0 56764 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_618
timestamp 1666464484
transform 1 0 57960 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_624
timestamp 1666464484
transform 1 0 58512 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1666464484
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1666464484
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1666464484
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1666464484
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_246
timestamp 1666464484
transform 1 0 23736 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_259
timestamp 1666464484
transform 1 0 24932 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_269
timestamp 1666464484
transform 1 0 25852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1666464484
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_289
timestamp 1666464484
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1666464484
transform 1 0 28152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_300
timestamp 1666464484
transform 1 0 28704 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_311
timestamp 1666464484
transform 1 0 29716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_325
timestamp 1666464484
transform 1 0 31004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1666464484
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_346
timestamp 1666464484
transform 1 0 32936 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_356
timestamp 1666464484
transform 1 0 33856 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_368
timestamp 1666464484
transform 1 0 34960 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_376
timestamp 1666464484
transform 1 0 35696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_382
timestamp 1666464484
transform 1 0 36248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1666464484
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_405
timestamp 1666464484
transform 1 0 38364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_415
timestamp 1666464484
transform 1 0 39284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_421
timestamp 1666464484
transform 1 0 39836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_435
timestamp 1666464484
transform 1 0 41124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_442
timestamp 1666464484
transform 1 0 41768 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_454
timestamp 1666464484
transform 1 0 42872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_460
timestamp 1666464484
transform 1 0 43424 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_468
timestamp 1666464484
transform 1 0 44160 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_476
timestamp 1666464484
transform 1 0 44896 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_489
timestamp 1666464484
transform 1 0 46092 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1666464484
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666464484
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_509
timestamp 1666464484
transform 1 0 47932 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_515
timestamp 1666464484
transform 1 0 48484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_525
timestamp 1666464484
transform 1 0 49404 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_531
timestamp 1666464484
transform 1 0 49956 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_536
timestamp 1666464484
transform 1 0 50416 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_550
timestamp 1666464484
transform 1 0 51704 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_556
timestamp 1666464484
transform 1 0 52256 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_561
timestamp 1666464484
transform 1 0 52716 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_567
timestamp 1666464484
transform 1 0 53268 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_575
timestamp 1666464484
transform 1 0 54004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_584
timestamp 1666464484
transform 1 0 54832 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_598
timestamp 1666464484
transform 1 0 56120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_602
timestamp 1666464484
transform 1 0 56488 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_606
timestamp 1666464484
transform 1 0 56856 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_612
timestamp 1666464484
transform 1 0 57408 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_617
timestamp 1666464484
transform 1 0 57868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_623
timestamp 1666464484
transform 1 0 58420 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1666464484
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1666464484
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1666464484
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1666464484
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1666464484
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1666464484
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_260
timestamp 1666464484
transform 1 0 25024 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_268
timestamp 1666464484
transform 1 0 25760 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_285
timestamp 1666464484
transform 1 0 27324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_293
timestamp 1666464484
transform 1 0 28060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1666464484
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666464484
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_318
timestamp 1666464484
transform 1 0 30360 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_326
timestamp 1666464484
transform 1 0 31096 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_334
timestamp 1666464484
transform 1 0 31832 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_341
timestamp 1666464484
transform 1 0 32476 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_345
timestamp 1666464484
transform 1 0 32844 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_351
timestamp 1666464484
transform 1 0 33396 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1666464484
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_371
timestamp 1666464484
transform 1 0 35236 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_379
timestamp 1666464484
transform 1 0 35972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_385
timestamp 1666464484
transform 1 0 36524 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_393
timestamp 1666464484
transform 1 0 37260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_397
timestamp 1666464484
transform 1 0 37628 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_408
timestamp 1666464484
transform 1 0 38640 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_433
timestamp 1666464484
transform 1 0 40940 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_437
timestamp 1666464484
transform 1 0 41308 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_440
timestamp 1666464484
transform 1 0 41584 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_450
timestamp 1666464484
transform 1 0 42504 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1666464484
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_477
timestamp 1666464484
transform 1 0 44988 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_481
timestamp 1666464484
transform 1 0 45356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_487
timestamp 1666464484
transform 1 0 45908 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_493
timestamp 1666464484
transform 1 0 46460 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_497
timestamp 1666464484
transform 1 0 46828 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_505
timestamp 1666464484
transform 1 0 47564 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_512
timestamp 1666464484
transform 1 0 48208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_516
timestamp 1666464484
transform 1 0 48576 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_523
timestamp 1666464484
transform 1 0 49220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_533
timestamp 1666464484
transform 1 0 50140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_549
timestamp 1666464484
transform 1 0 51612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_560
timestamp 1666464484
transform 1 0 52624 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_570
timestamp 1666464484
transform 1 0 53544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_580
timestamp 1666464484
transform 1 0 54464 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_589
timestamp 1666464484
transform 1 0 55292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_598
timestamp 1666464484
transform 1 0 56120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_607
timestamp 1666464484
transform 1 0 56948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_618
timestamp 1666464484
transform 1 0 57960 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_624
timestamp 1666464484
transform 1 0 58512 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1666464484
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1666464484
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1666464484
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1666464484
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1666464484
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1666464484
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1666464484
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1666464484
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_245
timestamp 1666464484
transform 1 0 23644 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_253
timestamp 1666464484
transform 1 0 24380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_260
timestamp 1666464484
transform 1 0 25024 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_267
timestamp 1666464484
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1666464484
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_285
timestamp 1666464484
transform 1 0 27324 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_296
timestamp 1666464484
transform 1 0 28336 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_308
timestamp 1666464484
transform 1 0 29440 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_322
timestamp 1666464484
transform 1 0 30728 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1666464484
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_343
timestamp 1666464484
transform 1 0 32660 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_349
timestamp 1666464484
transform 1 0 33212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_353
timestamp 1666464484
transform 1 0 33580 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_357
timestamp 1666464484
transform 1 0 33948 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_363
timestamp 1666464484
transform 1 0 34500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_371
timestamp 1666464484
transform 1 0 35236 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_377
timestamp 1666464484
transform 1 0 35788 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_383
timestamp 1666464484
transform 1 0 36340 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1666464484
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666464484
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_402
timestamp 1666464484
transform 1 0 38088 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_413
timestamp 1666464484
transform 1 0 39100 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_425
timestamp 1666464484
transform 1 0 40204 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_431
timestamp 1666464484
transform 1 0 40756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_438
timestamp 1666464484
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1666464484
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_464
timestamp 1666464484
transform 1 0 43792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_493
timestamp 1666464484
transform 1 0 46460 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_499
timestamp 1666464484
transform 1 0 47012 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666464484
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_510
timestamp 1666464484
transform 1 0 48024 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_525
timestamp 1666464484
transform 1 0 49404 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_537
timestamp 1666464484
transform 1 0 50508 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_549
timestamp 1666464484
transform 1 0 51612 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_557
timestamp 1666464484
transform 1 0 52348 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1666464484
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_573
timestamp 1666464484
transform 1 0 53820 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_582
timestamp 1666464484
transform 1 0 54648 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_589
timestamp 1666464484
transform 1 0 55292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_601
timestamp 1666464484
transform 1 0 56396 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_605
timestamp 1666464484
transform 1 0 56764 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1666464484
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1666464484
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_617
timestamp 1666464484
transform 1 0 57868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_622
timestamp 1666464484
transform 1 0 58328 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1666464484
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1666464484
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1666464484
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1666464484
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1666464484
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_245
timestamp 1666464484
transform 1 0 23644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1666464484
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_262
timestamp 1666464484
transform 1 0 25208 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_275
timestamp 1666464484
transform 1 0 26404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_281
timestamp 1666464484
transform 1 0 26956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1666464484
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_298
timestamp 1666464484
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1666464484
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_321
timestamp 1666464484
transform 1 0 30636 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_328
timestamp 1666464484
transform 1 0 31280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_340
timestamp 1666464484
transform 1 0 32384 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_348
timestamp 1666464484
transform 1 0 33120 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1666464484
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666464484
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1666464484
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_401
timestamp 1666464484
transform 1 0 37996 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_409
timestamp 1666464484
transform 1 0 38732 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_418
timestamp 1666464484
transform 1 0 39560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_427
timestamp 1666464484
transform 1 0 40388 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_436
timestamp 1666464484
transform 1 0 41216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_447
timestamp 1666464484
transform 1 0 42228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_451
timestamp 1666464484
transform 1 0 42596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_454
timestamp 1666464484
transform 1 0 42872 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_460
timestamp 1666464484
transform 1 0 43424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_463
timestamp 1666464484
transform 1 0 43700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_467
timestamp 1666464484
transform 1 0 44068 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1666464484
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_477
timestamp 1666464484
transform 1 0 44988 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_485
timestamp 1666464484
transform 1 0 45724 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_490
timestamp 1666464484
transform 1 0 46184 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_503
timestamp 1666464484
transform 1 0 47380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_515
timestamp 1666464484
transform 1 0 48484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_526
timestamp 1666464484
transform 1 0 49496 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_533
timestamp 1666464484
transform 1 0 50140 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_542
timestamp 1666464484
transform 1 0 50968 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_554
timestamp 1666464484
transform 1 0 52072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_563
timestamp 1666464484
transform 1 0 52900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_574
timestamp 1666464484
transform 1 0 53912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1666464484
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1666464484
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_589
timestamp 1666464484
transform 1 0 55292 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_596
timestamp 1666464484
transform 1 0 55936 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_606
timestamp 1666464484
transform 1 0 56856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_614
timestamp 1666464484
transform 1 0 57592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_622
timestamp 1666464484
transform 1 0 58328 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1666464484
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1666464484
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1666464484
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1666464484
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1666464484
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_237
timestamp 1666464484
transform 1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_245
timestamp 1666464484
transform 1 0 23644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_257
timestamp 1666464484
transform 1 0 24748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_261
timestamp 1666464484
transform 1 0 25116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1666464484
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_293
timestamp 1666464484
transform 1 0 28060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_297
timestamp 1666464484
transform 1 0 28428 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_304
timestamp 1666464484
transform 1 0 29072 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1666464484
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666464484
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_345
timestamp 1666464484
transform 1 0 32844 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_368
timestamp 1666464484
transform 1 0 34960 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_380
timestamp 1666464484
transform 1 0 36064 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_400
timestamp 1666464484
transform 1 0 37904 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_412
timestamp 1666464484
transform 1 0 39008 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_417
timestamp 1666464484
transform 1 0 39468 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_424
timestamp 1666464484
transform 1 0 40112 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_431
timestamp 1666464484
transform 1 0 40756 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_438
timestamp 1666464484
transform 1 0 41400 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1666464484
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_471
timestamp 1666464484
transform 1 0 44436 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_477
timestamp 1666464484
transform 1 0 44988 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_481
timestamp 1666464484
transform 1 0 45356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_490
timestamp 1666464484
transform 1 0 46184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_496
timestamp 1666464484
transform 1 0 46736 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_502
timestamp 1666464484
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_514
timestamp 1666464484
transform 1 0 48392 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_522
timestamp 1666464484
transform 1 0 49128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_527
timestamp 1666464484
transform 1 0 49588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_535
timestamp 1666464484
transform 1 0 50324 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_543
timestamp 1666464484
transform 1 0 51060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_547
timestamp 1666464484
transform 1 0 51428 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_555
timestamp 1666464484
transform 1 0 52164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1666464484
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_561
timestamp 1666464484
transform 1 0 52716 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_567
timestamp 1666464484
transform 1 0 53268 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_578
timestamp 1666464484
transform 1 0 54280 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_584
timestamp 1666464484
transform 1 0 54832 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_588
timestamp 1666464484
transform 1 0 55200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_598
timestamp 1666464484
transform 1 0 56120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_602
timestamp 1666464484
transform 1 0 56488 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_608
timestamp 1666464484
transform 1 0 57040 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_617
timestamp 1666464484
transform 1 0 57868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_621
timestamp 1666464484
transform 1 0 58236 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1666464484
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1666464484
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1666464484
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_233
timestamp 1666464484
transform 1 0 22540 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1666464484
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_265
timestamp 1666464484
transform 1 0 25484 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_293
timestamp 1666464484
transform 1 0 28060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1666464484
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666464484
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_317
timestamp 1666464484
transform 1 0 30268 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_321
timestamp 1666464484
transform 1 0 30636 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_327
timestamp 1666464484
transform 1 0 31188 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_338
timestamp 1666464484
transform 1 0 32200 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_350
timestamp 1666464484
transform 1 0 33304 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_358
timestamp 1666464484
transform 1 0 34040 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1666464484
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_373
timestamp 1666464484
transform 1 0 35420 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_379
timestamp 1666464484
transform 1 0 35972 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_387
timestamp 1666464484
transform 1 0 36708 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_398
timestamp 1666464484
transform 1 0 37720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_408
timestamp 1666464484
transform 1 0 38640 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_416
timestamp 1666464484
transform 1 0 39376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_437
timestamp 1666464484
transform 1 0 41308 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_461
timestamp 1666464484
transform 1 0 43516 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1666464484
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_477
timestamp 1666464484
transform 1 0 44988 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_485
timestamp 1666464484
transform 1 0 45724 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_494
timestamp 1666464484
transform 1 0 46552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_502
timestamp 1666464484
transform 1 0 47288 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_512
timestamp 1666464484
transform 1 0 48208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_516
timestamp 1666464484
transform 1 0 48576 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_521
timestamp 1666464484
transform 1 0 49036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_525
timestamp 1666464484
transform 1 0 49404 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_530
timestamp 1666464484
transform 1 0 49864 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_533
timestamp 1666464484
transform 1 0 50140 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_537
timestamp 1666464484
transform 1 0 50508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_549
timestamp 1666464484
transform 1 0 51612 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_557
timestamp 1666464484
transform 1 0 52348 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_565
timestamp 1666464484
transform 1 0 53084 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_573
timestamp 1666464484
transform 1 0 53820 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_585
timestamp 1666464484
transform 1 0 54924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_589
timestamp 1666464484
transform 1 0 55292 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_598
timestamp 1666464484
transform 1 0 56120 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_615
timestamp 1666464484
transform 1 0 57684 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_622
timestamp 1666464484
transform 1 0 58328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_9
timestamp 1666464484
transform 1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1666464484
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1666464484
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1666464484
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1666464484
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1666464484
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_249
timestamp 1666464484
transform 1 0 24012 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_268
timestamp 1666464484
transform 1 0 25760 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_302
timestamp 1666464484
transform 1 0 28888 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_319
timestamp 1666464484
transform 1 0 30452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_327
timestamp 1666464484
transform 1 0 31188 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1666464484
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1666464484
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_361
timestamp 1666464484
transform 1 0 34316 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_367
timestamp 1666464484
transform 1 0 34868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_372
timestamp 1666464484
transform 1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_379
timestamp 1666464484
transform 1 0 35972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_386
timestamp 1666464484
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_405
timestamp 1666464484
transform 1 0 38364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_414
timestamp 1666464484
transform 1 0 39192 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_429
timestamp 1666464484
transform 1 0 40572 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_436
timestamp 1666464484
transform 1 0 41216 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_442
timestamp 1666464484
transform 1 0 41768 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_454
timestamp 1666464484
transform 1 0 42872 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_462
timestamp 1666464484
transform 1 0 43608 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_467
timestamp 1666464484
transform 1 0 44068 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_475
timestamp 1666464484
transform 1 0 44804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_482
timestamp 1666464484
transform 1 0 45448 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_488
timestamp 1666464484
transform 1 0 46000 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_494
timestamp 1666464484
transform 1 0 46552 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_501
timestamp 1666464484
transform 1 0 47196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_512
timestamp 1666464484
transform 1 0 48208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_521
timestamp 1666464484
transform 1 0 49036 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_531
timestamp 1666464484
transform 1 0 49956 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_535
timestamp 1666464484
transform 1 0 50324 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_541
timestamp 1666464484
transform 1 0 50876 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_550
timestamp 1666464484
transform 1 0 51704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_558
timestamp 1666464484
transform 1 0 52440 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_561
timestamp 1666464484
transform 1 0 52716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_567
timestamp 1666464484
transform 1 0 53268 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_578
timestamp 1666464484
transform 1 0 54280 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_590
timestamp 1666464484
transform 1 0 55384 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_598
timestamp 1666464484
transform 1 0 56120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_603
timestamp 1666464484
transform 1 0 56580 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_607
timestamp 1666464484
transform 1 0 56948 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_614
timestamp 1666464484
transform 1 0 57592 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_617
timestamp 1666464484
transform 1 0 57868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_623
timestamp 1666464484
transform 1 0 58420 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1666464484
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1666464484
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1666464484
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1666464484
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666464484
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666464484
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1666464484
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_285
timestamp 1666464484
transform 1 0 27324 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_290
timestamp 1666464484
transform 1 0 27784 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1666464484
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_321
timestamp 1666464484
transform 1 0 30636 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_327
timestamp 1666464484
transform 1 0 31188 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_350
timestamp 1666464484
transform 1 0 33304 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1666464484
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_376
timestamp 1666464484
transform 1 0 35696 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_384
timestamp 1666464484
transform 1 0 36432 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_392
timestamp 1666464484
transform 1 0 37168 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_404
timestamp 1666464484
transform 1 0 38272 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_408
timestamp 1666464484
transform 1 0 38640 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_431
timestamp 1666464484
transform 1 0 40756 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_443
timestamp 1666464484
transform 1 0 41860 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_455
timestamp 1666464484
transform 1 0 42964 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_460
timestamp 1666464484
transform 1 0 43424 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_468
timestamp 1666464484
transform 1 0 44160 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1666464484
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_484
timestamp 1666464484
transform 1 0 45632 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_492
timestamp 1666464484
transform 1 0 46368 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_498
timestamp 1666464484
transform 1 0 46920 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_504
timestamp 1666464484
transform 1 0 47472 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_507
timestamp 1666464484
transform 1 0 47748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_519
timestamp 1666464484
transform 1 0 48852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_533
timestamp 1666464484
transform 1 0 50140 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_543
timestamp 1666464484
transform 1 0 51060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_555
timestamp 1666464484
transform 1 0 52164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_563
timestamp 1666464484
transform 1 0 52900 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_571
timestamp 1666464484
transform 1 0 53636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_586
timestamp 1666464484
transform 1 0 55016 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_589
timestamp 1666464484
transform 1 0 55292 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_596
timestamp 1666464484
transform 1 0 55936 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_610
timestamp 1666464484
transform 1 0 57224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_620
timestamp 1666464484
transform 1 0 58144 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_624
timestamp 1666464484
transform 1 0 58512 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666464484
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1666464484
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1666464484
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1666464484
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666464484
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1666464484
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1666464484
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1666464484
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1666464484
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1666464484
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_361
timestamp 1666464484
transform 1 0 34316 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_373
timestamp 1666464484
transform 1 0 35420 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_377
timestamp 1666464484
transform 1 0 35788 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1666464484
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666464484
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_400
timestamp 1666464484
transform 1 0 37904 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_412
timestamp 1666464484
transform 1 0 39008 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_427
timestamp 1666464484
transform 1 0 40388 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_439
timestamp 1666464484
transform 1 0 41492 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666464484
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_465
timestamp 1666464484
transform 1 0 43884 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_476
timestamp 1666464484
transform 1 0 44896 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_480
timestamp 1666464484
transform 1 0 45264 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_488
timestamp 1666464484
transform 1 0 46000 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_496
timestamp 1666464484
transform 1 0 46736 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_502
timestamp 1666464484
transform 1 0 47288 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_512
timestamp 1666464484
transform 1 0 48208 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_523
timestamp 1666464484
transform 1 0 49220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_538
timestamp 1666464484
transform 1 0 50600 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_550
timestamp 1666464484
transform 1 0 51704 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_554
timestamp 1666464484
transform 1 0 52072 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_558
timestamp 1666464484
transform 1 0 52440 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_561
timestamp 1666464484
transform 1 0 52716 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_569
timestamp 1666464484
transform 1 0 53452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_581
timestamp 1666464484
transform 1 0 54556 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_604
timestamp 1666464484
transform 1 0 56672 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_611
timestamp 1666464484
transform 1 0 57316 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1666464484
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_617
timestamp 1666464484
transform 1 0 57868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1666464484
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1666464484
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1666464484
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1666464484
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1666464484
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1666464484
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1666464484
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1666464484
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666464484
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1666464484
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1666464484
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1666464484
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1666464484
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1666464484
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666464484
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_389
timestamp 1666464484
transform 1 0 36892 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_396
timestamp 1666464484
transform 1 0 37536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_400
timestamp 1666464484
transform 1 0 37904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_406
timestamp 1666464484
transform 1 0 38456 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_417
timestamp 1666464484
transform 1 0 39468 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_428
timestamp 1666464484
transform 1 0 40480 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_440
timestamp 1666464484
transform 1 0 41584 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_452
timestamp 1666464484
transform 1 0 42688 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_460
timestamp 1666464484
transform 1 0 43424 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_466
timestamp 1666464484
transform 1 0 43976 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_472
timestamp 1666464484
transform 1 0 44528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_477
timestamp 1666464484
transform 1 0 44988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_486
timestamp 1666464484
transform 1 0 45816 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_492
timestamp 1666464484
transform 1 0 46368 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_498
timestamp 1666464484
transform 1 0 46920 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_506
timestamp 1666464484
transform 1 0 47656 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_512
timestamp 1666464484
transform 1 0 48208 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_520
timestamp 1666464484
transform 1 0 48944 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_530
timestamp 1666464484
transform 1 0 49864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_533
timestamp 1666464484
transform 1 0 50140 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_542
timestamp 1666464484
transform 1 0 50968 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_567
timestamp 1666464484
transform 1 0 53268 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_573
timestamp 1666464484
transform 1 0 53820 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_577
timestamp 1666464484
transform 1 0 54188 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_585
timestamp 1666464484
transform 1 0 54924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_589
timestamp 1666464484
transform 1 0 55292 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_599
timestamp 1666464484
transform 1 0 56212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_603
timestamp 1666464484
transform 1 0 56580 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_606
timestamp 1666464484
transform 1 0 56856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_623
timestamp 1666464484
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1666464484
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1666464484
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1666464484
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1666464484
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1666464484
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1666464484
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1666464484
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666464484
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666464484
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666464484
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666464484
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_401
timestamp 1666464484
transform 1 0 37996 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_424
timestamp 1666464484
transform 1 0 40112 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_436
timestamp 1666464484
transform 1 0 41216 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_474
timestamp 1666464484
transform 1 0 44712 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_481
timestamp 1666464484
transform 1 0 45356 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_490
timestamp 1666464484
transform 1 0 46184 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_498
timestamp 1666464484
transform 1 0 46920 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_509
timestamp 1666464484
transform 1 0 47932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_515
timestamp 1666464484
transform 1 0 48484 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_521
timestamp 1666464484
transform 1 0 49036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_544
timestamp 1666464484
transform 1 0 51152 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_556
timestamp 1666464484
transform 1 0 52256 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_561
timestamp 1666464484
transform 1 0 52716 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_568
timestamp 1666464484
transform 1 0 53360 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_579
timestamp 1666464484
transform 1 0 54372 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_588
timestamp 1666464484
transform 1 0 55200 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_596
timestamp 1666464484
transform 1 0 55936 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_602
timestamp 1666464484
transform 1 0 56488 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_614
timestamp 1666464484
transform 1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_617
timestamp 1666464484
transform 1 0 57868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_622
timestamp 1666464484
transform 1 0 58328 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1666464484
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1666464484
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1666464484
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1666464484
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1666464484
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1666464484
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1666464484
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666464484
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666464484
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666464484
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1666464484
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1666464484
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666464484
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666464484
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666464484
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_401
timestamp 1666464484
transform 1 0 37996 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_405
timestamp 1666464484
transform 1 0 38364 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_412
timestamp 1666464484
transform 1 0 39008 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666464484
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666464484
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_457
timestamp 1666464484
transform 1 0 43148 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_465
timestamp 1666464484
transform 1 0 43884 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_472
timestamp 1666464484
transform 1 0 44528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_477
timestamp 1666464484
transform 1 0 44988 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_485
timestamp 1666464484
transform 1 0 45724 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_494
timestamp 1666464484
transform 1 0 46552 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_503
timestamp 1666464484
transform 1 0 47380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_512
timestamp 1666464484
transform 1 0 48208 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_528
timestamp 1666464484
transform 1 0 49680 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_533
timestamp 1666464484
transform 1 0 50140 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_537
timestamp 1666464484
transform 1 0 50508 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_542
timestamp 1666464484
transform 1 0 50968 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_554
timestamp 1666464484
transform 1 0 52072 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_562
timestamp 1666464484
transform 1 0 52808 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_586
timestamp 1666464484
transform 1 0 55016 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_589
timestamp 1666464484
transform 1 0 55292 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_613
timestamp 1666464484
transform 1 0 57500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_622
timestamp 1666464484
transform 1 0 58328 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1666464484
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1666464484
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1666464484
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666464484
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666464484
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1666464484
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1666464484
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1666464484
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1666464484
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666464484
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666464484
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666464484
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1666464484
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666464484
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666464484
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666464484
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666464484
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666464484
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_457
timestamp 1666464484
transform 1 0 43148 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_464
timestamp 1666464484
transform 1 0 43792 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_483
timestamp 1666464484
transform 1 0 45540 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_491
timestamp 1666464484
transform 1 0 46276 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666464484
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666464484
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_514
timestamp 1666464484
transform 1 0 48392 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_526
timestamp 1666464484
transform 1 0 49496 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_531
timestamp 1666464484
transform 1 0 49956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_539
timestamp 1666464484
transform 1 0 50692 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_545
timestamp 1666464484
transform 1 0 51244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_558
timestamp 1666464484
transform 1 0 52440 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_561
timestamp 1666464484
transform 1 0 52716 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_569
timestamp 1666464484
transform 1 0 53452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_577
timestamp 1666464484
transform 1 0 54188 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_581
timestamp 1666464484
transform 1 0 54556 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_587
timestamp 1666464484
transform 1 0 55108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_591
timestamp 1666464484
transform 1 0 55476 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_598
timestamp 1666464484
transform 1 0 56120 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_606
timestamp 1666464484
transform 1 0 56856 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_614
timestamp 1666464484
transform 1 0 57592 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1666464484
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1666464484
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666464484
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666464484
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1666464484
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666464484
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1666464484
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1666464484
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1666464484
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1666464484
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666464484
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666464484
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666464484
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666464484
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666464484
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666464484
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666464484
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666464484
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_457
timestamp 1666464484
transform 1 0 43148 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_474
timestamp 1666464484
transform 1 0 44712 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_477
timestamp 1666464484
transform 1 0 44988 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_490
timestamp 1666464484
transform 1 0 46184 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_496
timestamp 1666464484
transform 1 0 46736 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_502
timestamp 1666464484
transform 1 0 47288 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_513
timestamp 1666464484
transform 1 0 48300 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_521
timestamp 1666464484
transform 1 0 49036 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_529
timestamp 1666464484
transform 1 0 49772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_533
timestamp 1666464484
transform 1 0 50140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_537
timestamp 1666464484
transform 1 0 50508 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_544
timestamp 1666464484
transform 1 0 51152 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_565
timestamp 1666464484
transform 1 0 53084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_569
timestamp 1666464484
transform 1 0 53452 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_577
timestamp 1666464484
transform 1 0 54188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_584
timestamp 1666464484
transform 1 0 54832 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_589
timestamp 1666464484
transform 1 0 55292 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_594
timestamp 1666464484
transform 1 0 55752 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_600
timestamp 1666464484
transform 1 0 56304 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_623
timestamp 1666464484
transform 1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1666464484
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666464484
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666464484
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666464484
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666464484
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666464484
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666464484
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666464484
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666464484
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1666464484
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1666464484
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1666464484
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1666464484
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666464484
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666464484
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666464484
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666464484
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666464484
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666464484
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666464484
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666464484
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666464484
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_461
timestamp 1666464484
transform 1 0 43516 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_484
timestamp 1666464484
transform 1 0 45632 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_495
timestamp 1666464484
transform 1 0 46644 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_501
timestamp 1666464484
transform 1 0 47196 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_516
timestamp 1666464484
transform 1 0 48576 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_538
timestamp 1666464484
transform 1 0 50600 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_549
timestamp 1666464484
transform 1 0 51612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_558
timestamp 1666464484
transform 1 0 52440 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_561
timestamp 1666464484
transform 1 0 52716 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_584
timestamp 1666464484
transform 1 0 54832 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_610
timestamp 1666464484
transform 1 0 57224 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1666464484
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666464484
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666464484
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1666464484
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666464484
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666464484
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666464484
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1666464484
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666464484
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666464484
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666464484
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666464484
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666464484
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666464484
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666464484
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666464484
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666464484
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666464484
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666464484
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666464484
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666464484
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666464484
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666464484
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666464484
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_477
timestamp 1666464484
transform 1 0 44988 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_485
timestamp 1666464484
transform 1 0 45724 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_492
timestamp 1666464484
transform 1 0 46368 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_502
timestamp 1666464484
transform 1 0 47288 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_514
timestamp 1666464484
transform 1 0 48392 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_522
timestamp 1666464484
transform 1 0 49128 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_530
timestamp 1666464484
transform 1 0 49864 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_533
timestamp 1666464484
transform 1 0 50140 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_540
timestamp 1666464484
transform 1 0 50784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_565
timestamp 1666464484
transform 1 0 53084 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_569
timestamp 1666464484
transform 1 0 53452 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_575
timestamp 1666464484
transform 1 0 54004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1666464484
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1666464484
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_601
timestamp 1666464484
transform 1 0 56396 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_608
timestamp 1666464484
transform 1 0 57040 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_620
timestamp 1666464484
transform 1 0 58144 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_624
timestamp 1666464484
transform 1 0 58512 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1666464484
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1666464484
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666464484
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1666464484
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1666464484
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1666464484
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666464484
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666464484
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1666464484
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1666464484
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1666464484
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666464484
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666464484
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666464484
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666464484
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666464484
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666464484
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666464484
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666464484
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666464484
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666464484
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666464484
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666464484
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_461
timestamp 1666464484
transform 1 0 43516 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_467
timestamp 1666464484
transform 1 0 44068 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_481
timestamp 1666464484
transform 1 0 45356 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_492
timestamp 1666464484
transform 1 0 46368 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_502
timestamp 1666464484
transform 1 0 47288 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_515
timestamp 1666464484
transform 1 0 48484 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_521
timestamp 1666464484
transform 1 0 49036 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_543
timestamp 1666464484
transform 1 0 51060 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_552
timestamp 1666464484
transform 1 0 51888 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_561
timestamp 1666464484
transform 1 0 52716 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_586
timestamp 1666464484
transform 1 0 55016 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_598
timestamp 1666464484
transform 1 0 56120 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_610
timestamp 1666464484
transform 1 0 57224 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1666464484
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_9
timestamp 1666464484
transform 1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1666464484
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1666464484
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1666464484
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1666464484
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1666464484
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1666464484
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666464484
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666464484
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666464484
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666464484
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666464484
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666464484
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1666464484
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1666464484
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1666464484
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1666464484
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666464484
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666464484
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1666464484
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1666464484
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666464484
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_477
timestamp 1666464484
transform 1 0 44988 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_487
timestamp 1666464484
transform 1 0 45908 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_497
timestamp 1666464484
transform 1 0 46828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_504
timestamp 1666464484
transform 1 0 47472 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_514
timestamp 1666464484
transform 1 0 48392 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_524
timestamp 1666464484
transform 1 0 49312 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_533
timestamp 1666464484
transform 1 0 50140 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_539
timestamp 1666464484
transform 1 0 50692 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_543
timestamp 1666464484
transform 1 0 51060 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_554
timestamp 1666464484
transform 1 0 52072 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_566
timestamp 1666464484
transform 1 0 53176 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_578
timestamp 1666464484
transform 1 0 54280 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_586
timestamp 1666464484
transform 1 0 55016 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1666464484
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1666464484
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1666464484
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1666464484
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1666464484
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1666464484
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1666464484
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666464484
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666464484
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666464484
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666464484
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666464484
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666464484
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666464484
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1666464484
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1666464484
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1666464484
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1666464484
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666464484
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666464484
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_473
timestamp 1666464484
transform 1 0 44620 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_481
timestamp 1666464484
transform 1 0 45356 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_496
timestamp 1666464484
transform 1 0 46736 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_517
timestamp 1666464484
transform 1 0 48668 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_530
timestamp 1666464484
transform 1 0 49864 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_542
timestamp 1666464484
transform 1 0 50968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_554
timestamp 1666464484
transform 1 0 52072 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1666464484
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1666464484
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1666464484
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1666464484
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1666464484
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1666464484
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1666464484
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1666464484
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1666464484
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1666464484
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1666464484
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1666464484
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666464484
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1666464484
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1666464484
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1666464484
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1666464484
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1666464484
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1666464484
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1666464484
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666464484
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1666464484
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1666464484
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1666464484
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1666464484
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666464484
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666464484
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666464484
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666464484
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666464484
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_477
timestamp 1666464484
transform 1 0 44988 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_507
timestamp 1666464484
transform 1 0 47748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_524
timestamp 1666464484
transform 1 0 49312 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1666464484
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1666464484
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1666464484
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1666464484
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1666464484
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1666464484
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1666464484
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1666464484
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_613
timestamp 1666464484
transform 1 0 57500 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_623
timestamp 1666464484
transform 1 0 58420 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1666464484
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1666464484
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666464484
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666464484
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1666464484
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1666464484
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1666464484
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1666464484
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1666464484
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1666464484
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1666464484
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1666464484
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666464484
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666464484
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666464484
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666464484
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1666464484
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1666464484
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1666464484
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1666464484
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666464484
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666464484
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666464484
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666464484
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666464484
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666464484
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_461
timestamp 1666464484
transform 1 0 43516 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_491
timestamp 1666464484
transform 1 0 46276 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_500
timestamp 1666464484
transform 1 0 47104 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1666464484
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1666464484
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1666464484
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1666464484
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1666464484
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1666464484
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1666464484
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1666464484
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1666464484
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666464484
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1666464484
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1666464484
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1666464484
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1666464484
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1666464484
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666464484
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1666464484
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1666464484
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1666464484
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1666464484
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666464484
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666464484
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666464484
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666464484
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666464484
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666464484
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666464484
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1666464484
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1666464484
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1666464484
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666464484
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666464484
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666464484
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666464484
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1666464484
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1666464484
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1666464484
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1666464484
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1666464484
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1666464484
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1666464484
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1666464484
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1666464484
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1666464484
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1666464484
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1666464484
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1666464484
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1666464484
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1666464484
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1666464484
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666464484
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1666464484
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1666464484
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1666464484
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1666464484
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666464484
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666464484
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666464484
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1666464484
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666464484
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666464484
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1666464484
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1666464484
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1666464484
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1666464484
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666464484
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666464484
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666464484
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666464484
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666464484
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666464484
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666464484
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1666464484
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1666464484
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1666464484
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666464484
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1666464484
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1666464484
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1666464484
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1666464484
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1666464484
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1666464484
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1666464484
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1666464484
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1666464484
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1666464484
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1666464484
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1666464484
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1666464484
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1666464484
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666464484
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666464484
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666464484
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1666464484
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1666464484
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666464484
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666464484
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666464484
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666464484
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666464484
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666464484
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666464484
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1666464484
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1666464484
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1666464484
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666464484
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666464484
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666464484
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666464484
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1666464484
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1666464484
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1666464484
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1666464484
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1666464484
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1666464484
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1666464484
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1666464484
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1666464484
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1666464484
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1666464484
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1666464484
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1666464484
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1666464484
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666464484
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1666464484
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1666464484
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1666464484
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1666464484
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666464484
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1666464484
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1666464484
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1666464484
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1666464484
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666464484
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1666464484
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1666464484
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1666464484
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1666464484
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666464484
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1666464484
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1666464484
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1666464484
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1666464484
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666464484
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666464484
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666464484
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666464484
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666464484
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666464484
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666464484
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666464484
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666464484
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666464484
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1666464484
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1666464484
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1666464484
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1666464484
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1666464484
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1666464484
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1666464484
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1666464484
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1666464484
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666464484
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1666464484
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1666464484
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666464484
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1666464484
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1666464484
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1666464484
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1666464484
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666464484
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1666464484
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1666464484
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1666464484
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1666464484
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666464484
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666464484
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1666464484
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1666464484
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1666464484
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666464484
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666464484
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666464484
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666464484
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666464484
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666464484
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1666464484
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1666464484
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1666464484
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1666464484
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666464484
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666464484
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666464484
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666464484
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1666464484
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1666464484
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1666464484
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1666464484
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1666464484
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1666464484
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1666464484
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1666464484
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1666464484
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1666464484
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1666464484
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1666464484
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666464484
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666464484
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666464484
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666464484
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1666464484
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666464484
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1666464484
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1666464484
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666464484
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1666464484
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666464484
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666464484
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1666464484
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1666464484
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1666464484
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666464484
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1666464484
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666464484
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666464484
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1666464484
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666464484
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666464484
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666464484
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666464484
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666464484
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666464484
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666464484
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666464484
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666464484
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666464484
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1666464484
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1666464484
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1666464484
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1666464484
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1666464484
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1666464484
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1666464484
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1666464484
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1666464484
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1666464484
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1666464484
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666464484
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666464484
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1666464484
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1666464484
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1666464484
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1666464484
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666464484
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1666464484
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1666464484
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1666464484
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1666464484
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666464484
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1666464484
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1666464484
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1666464484
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1666464484
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666464484
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666464484
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666464484
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1666464484
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1666464484
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666464484
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1666464484
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1666464484
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1666464484
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1666464484
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666464484
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666464484
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666464484
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666464484
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666464484
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666464484
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666464484
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666464484
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666464484
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1666464484
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1666464484
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1666464484
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1666464484
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1666464484
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1666464484
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1666464484
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1666464484
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1666464484
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1666464484
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1666464484
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1666464484
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1666464484
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1666464484
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1666464484
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1666464484
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666464484
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666464484
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666464484
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1666464484
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1666464484
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666464484
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1666464484
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1666464484
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1666464484
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1666464484
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1666464484
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1666464484
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1666464484
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1666464484
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1666464484
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666464484
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1666464484
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1666464484
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1666464484
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1666464484
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666464484
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666464484
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666464484
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666464484
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666464484
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666464484
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666464484
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666464484
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666464484
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666464484
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1666464484
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1666464484
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1666464484
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1666464484
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1666464484
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1666464484
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1666464484
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1666464484
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1666464484
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1666464484
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1666464484
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1666464484
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666464484
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666464484
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666464484
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666464484
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1666464484
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1666464484
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666464484
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1666464484
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1666464484
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1666464484
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1666464484
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666464484
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1666464484
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1666464484
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1666464484
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1666464484
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666464484
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1666464484
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1666464484
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1666464484
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1666464484
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666464484
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666464484
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1666464484
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1666464484
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1666464484
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666464484
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666464484
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666464484
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666464484
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666464484
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666464484
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666464484
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666464484
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666464484
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1666464484
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1666464484
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1666464484
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1666464484
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1666464484
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1666464484
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1666464484
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1666464484
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1666464484
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1666464484
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1666464484
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1666464484
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1666464484
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1666464484
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666464484
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666464484
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666464484
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666464484
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666464484
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666464484
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666464484
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666464484
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666464484
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666464484
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1666464484
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1666464484
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666464484
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1666464484
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1666464484
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1666464484
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1666464484
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1666464484
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1666464484
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1666464484
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1666464484
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1666464484
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1666464484
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1666464484
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666464484
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666464484
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1666464484
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666464484
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666464484
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666464484
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666464484
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666464484
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666464484
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666464484
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1666464484
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1666464484
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1666464484
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666464484
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1666464484
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1666464484
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1666464484
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1666464484
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1666464484
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1666464484
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1666464484
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1666464484
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1666464484
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1666464484
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1666464484
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1666464484
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666464484
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666464484
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666464484
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666464484
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666464484
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666464484
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666464484
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666464484
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666464484
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666464484
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666464484
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666464484
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666464484
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666464484
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666464484
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1666464484
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1666464484
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1666464484
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1666464484
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666464484
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1666464484
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1666464484
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1666464484
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1666464484
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666464484
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1666464484
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1666464484
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1666464484
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1666464484
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666464484
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1666464484
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1666464484
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1666464484
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1666464484
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666464484
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666464484
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666464484
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666464484
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666464484
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666464484
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1666464484
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1666464484
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1666464484
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1666464484
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1666464484
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1666464484
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1666464484
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1666464484
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1666464484
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1666464484
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1666464484
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1666464484
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1666464484
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1666464484
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_613
timestamp 1666464484
transform 1 0 57500 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_64_623
timestamp 1666464484
transform 1 0 58420 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1666464484
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1666464484
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1666464484
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1666464484
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1666464484
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666464484
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666464484
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666464484
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666464484
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666464484
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666464484
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1666464484
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1666464484
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1666464484
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1666464484
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1666464484
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666464484
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666464484
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1666464484
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1666464484
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1666464484
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1666464484
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666464484
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1666464484
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1666464484
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1666464484
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1666464484
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1666464484
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666464484
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1666464484
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1666464484
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1666464484
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1666464484
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1666464484
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666464484
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1666464484
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1666464484
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1666464484
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1666464484
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1666464484
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666464484
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666464484
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666464484
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666464484
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666464484
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666464484
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666464484
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666464484
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666464484
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666464484
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666464484
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666464484
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666464484
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1666464484
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1666464484
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1666464484
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1666464484
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1666464484
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1666464484
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1666464484
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1666464484
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1666464484
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1666464484
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1666464484
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1666464484
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1666464484
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1666464484
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666464484
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666464484
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666464484
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666464484
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666464484
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666464484
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666464484
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666464484
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666464484
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666464484
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666464484
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666464484
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666464484
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666464484
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666464484
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666464484
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1666464484
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1666464484
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666464484
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1666464484
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1666464484
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1666464484
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1666464484
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1666464484
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1666464484
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1666464484
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1666464484
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1666464484
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1666464484
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1666464484
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1666464484
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1666464484
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1666464484
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1666464484
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1666464484
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1666464484
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666464484
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666464484
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1666464484
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1666464484
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666464484
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1666464484
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666464484
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666464484
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666464484
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666464484
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666464484
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666464484
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666464484
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666464484
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666464484
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666464484
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1666464484
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1666464484
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1666464484
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1666464484
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1666464484
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1666464484
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1666464484
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1666464484
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1666464484
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1666464484
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1666464484
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1666464484
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1666464484
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1666464484
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1666464484
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1666464484
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666464484
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666464484
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666464484
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666464484
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666464484
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666464484
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666464484
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666464484
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666464484
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1666464484
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1666464484
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1666464484
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666464484
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666464484
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1666464484
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1666464484
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666464484
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1666464484
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1666464484
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1666464484
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1666464484
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1666464484
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1666464484
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1666464484
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1666464484
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1666464484
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1666464484
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1666464484
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666464484
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1666464484
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1666464484
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666464484
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666464484
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1666464484
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1666464484
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666464484
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666464484
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666464484
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666464484
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666464484
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666464484
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666464484
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666464484
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666464484
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666464484
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666464484
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666464484
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1666464484
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1666464484
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1666464484
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1666464484
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1666464484
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1666464484
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1666464484
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1666464484
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1666464484
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1666464484
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1666464484
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1666464484
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1666464484
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1666464484
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666464484
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666464484
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666464484
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666464484
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666464484
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666464484
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666464484
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666464484
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666464484
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666464484
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666464484
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666464484
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666464484
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666464484
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666464484
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1666464484
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1666464484
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1666464484
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666464484
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666464484
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666464484
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1666464484
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1666464484
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1666464484
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666464484
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1666464484
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1666464484
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1666464484
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1666464484
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666464484
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666464484
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1666464484
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1666464484
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1666464484
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1666464484
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1666464484
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666464484
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1666464484
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666464484
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1666464484
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1666464484
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1666464484
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666464484
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666464484
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666464484
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666464484
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666464484
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666464484
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666464484
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666464484
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666464484
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666464484
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1666464484
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1666464484
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1666464484
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1666464484
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1666464484
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1666464484
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1666464484
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1666464484
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1666464484
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1666464484
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1666464484
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1666464484
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1666464484
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1666464484
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1666464484
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666464484
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666464484
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666464484
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666464484
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666464484
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666464484
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666464484
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666464484
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666464484
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666464484
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666464484
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666464484
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666464484
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666464484
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666464484
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666464484
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666464484
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666464484
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666464484
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1666464484
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1666464484
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1666464484
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1666464484
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1666464484
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1666464484
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1666464484
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1666464484
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1666464484
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1666464484
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1666464484
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666464484
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1666464484
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1666464484
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666464484
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666464484
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1666464484
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666464484
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666464484
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666464484
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666464484
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666464484
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666464484
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666464484
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666464484
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666464484
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666464484
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666464484
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666464484
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666464484
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1666464484
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1666464484
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1666464484
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1666464484
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1666464484
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1666464484
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1666464484
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1666464484
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1666464484
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1666464484
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1666464484
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1666464484
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1666464484
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1666464484
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666464484
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666464484
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666464484
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666464484
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666464484
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666464484
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666464484
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666464484
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666464484
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666464484
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666464484
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666464484
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666464484
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666464484
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666464484
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666464484
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1666464484
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1666464484
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666464484
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666464484
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666464484
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1666464484
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1666464484
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1666464484
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1666464484
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1666464484
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1666464484
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1666464484
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1666464484
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1666464484
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666464484
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1666464484
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1666464484
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1666464484
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1666464484
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1666464484
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666464484
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1666464484
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1666464484
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1666464484
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1666464484
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1666464484
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666464484
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666464484
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666464484
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666464484
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666464484
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666464484
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666464484
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666464484
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666464484
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666464484
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1666464484
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1666464484
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1666464484
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1666464484
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1666464484
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1666464484
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1666464484
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1666464484
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1666464484
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1666464484
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1666464484
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1666464484
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_9
timestamp 1666464484
transform 1 0 1932 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1666464484
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1666464484
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1666464484
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666464484
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666464484
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666464484
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666464484
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666464484
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666464484
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666464484
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666464484
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666464484
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666464484
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666464484
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666464484
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666464484
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666464484
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666464484
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666464484
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666464484
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1666464484
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666464484
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1666464484
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1666464484
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1666464484
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1666464484
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1666464484
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1666464484
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1666464484
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1666464484
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1666464484
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1666464484
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1666464484
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1666464484
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1666464484
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1666464484
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1666464484
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1666464484
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1666464484
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666464484
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666464484
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666464484
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666464484
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666464484
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666464484
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666464484
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666464484
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666464484
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666464484
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666464484
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666464484
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666464484
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1666464484
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1666464484
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1666464484
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1666464484
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1666464484
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1666464484
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1666464484
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1666464484
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1666464484
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1666464484
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1666464484
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1666464484
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1666464484
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1666464484
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666464484
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666464484
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666464484
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666464484
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666464484
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666464484
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666464484
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666464484
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666464484
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666464484
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666464484
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666464484
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666464484
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666464484
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666464484
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666464484
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666464484
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666464484
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666464484
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666464484
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1666464484
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1666464484
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1666464484
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1666464484
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1666464484
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1666464484
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1666464484
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1666464484
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1666464484
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1666464484
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1666464484
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1666464484
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1666464484
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1666464484
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1666464484
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1666464484
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1666464484
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1666464484
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1666464484
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1666464484
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1666464484
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1666464484
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1666464484
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666464484
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666464484
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666464484
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666464484
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666464484
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666464484
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666464484
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666464484
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666464484
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1666464484
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1666464484
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1666464484
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1666464484
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1666464484
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1666464484
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1666464484
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1666464484
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1666464484
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1666464484
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1666464484
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1666464484
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1666464484
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1666464484
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1666464484
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666464484
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666464484
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666464484
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666464484
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666464484
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666464484
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666464484
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666464484
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666464484
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666464484
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666464484
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666464484
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666464484
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666464484
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666464484
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666464484
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666464484
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1666464484
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666464484
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1666464484
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1666464484
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1666464484
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1666464484
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1666464484
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1666464484
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1666464484
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1666464484
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1666464484
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1666464484
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1666464484
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1666464484
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1666464484
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1666464484
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1666464484
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1666464484
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1666464484
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1666464484
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1666464484
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1666464484
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1666464484
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1666464484
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1666464484
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666464484
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666464484
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666464484
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666464484
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666464484
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666464484
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666464484
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1666464484
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1666464484
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1666464484
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1666464484
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1666464484
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1666464484
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1666464484
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1666464484
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1666464484
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1666464484
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1666464484
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1666464484
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1666464484
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1666464484
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666464484
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666464484
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666464484
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666464484
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666464484
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666464484
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666464484
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666464484
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666464484
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666464484
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666464484
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666464484
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666464484
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666464484
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666464484
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666464484
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666464484
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666464484
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666464484
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666464484
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666464484
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1666464484
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1666464484
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1666464484
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1666464484
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1666464484
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1666464484
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1666464484
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1666464484
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1666464484
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1666464484
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1666464484
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1666464484
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1666464484
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1666464484
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1666464484
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1666464484
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1666464484
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1666464484
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1666464484
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1666464484
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1666464484
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1666464484
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666464484
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666464484
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666464484
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666464484
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666464484
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666464484
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666464484
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666464484
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666464484
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1666464484
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1666464484
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1666464484
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1666464484
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1666464484
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1666464484
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1666464484
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1666464484
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1666464484
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1666464484
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1666464484
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_615
timestamp 1666464484
transform 1 0 57684 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_623
timestamp 1666464484
transform 1 0 58420 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1666464484
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1666464484
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1666464484
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1666464484
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1666464484
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666464484
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666464484
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666464484
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666464484
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666464484
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666464484
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666464484
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666464484
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666464484
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666464484
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666464484
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666464484
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666464484
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666464484
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666464484
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1666464484
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1666464484
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666464484
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1666464484
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1666464484
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1666464484
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1666464484
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1666464484
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1666464484
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1666464484
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1666464484
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1666464484
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1666464484
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1666464484
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1666464484
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1666464484
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1666464484
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1666464484
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1666464484
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1666464484
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1666464484
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1666464484
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1666464484
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1666464484
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1666464484
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1666464484
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1666464484
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666464484
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666464484
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666464484
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666464484
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666464484
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666464484
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1666464484
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1666464484
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1666464484
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1666464484
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1666464484
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1666464484
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1666464484
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1666464484
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1666464484
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1666464484
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1666464484
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1666464484
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666464484
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666464484
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666464484
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666464484
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666464484
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666464484
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666464484
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666464484
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666464484
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666464484
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666464484
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666464484
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666464484
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1666464484
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1666464484
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666464484
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666464484
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666464484
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666464484
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1666464484
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1666464484
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1666464484
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1666464484
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1666464484
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1666464484
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1666464484
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1666464484
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1666464484
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1666464484
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1666464484
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1666464484
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1666464484
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1666464484
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1666464484
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1666464484
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1666464484
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1666464484
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1666464484
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1666464484
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1666464484
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1666464484
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1666464484
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1666464484
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1666464484
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1666464484
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1666464484
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1666464484
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1666464484
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666464484
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666464484
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666464484
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666464484
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1666464484
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1666464484
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1666464484
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1666464484
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1666464484
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1666464484
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1666464484
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1666464484
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1666464484
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1666464484
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1666464484
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1666464484
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1666464484
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1666464484
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1666464484
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1666464484
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1666464484
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666464484
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666464484
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666464484
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666464484
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666464484
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666464484
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666464484
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666464484
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666464484
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666464484
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666464484
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666464484
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666464484
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666464484
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1666464484
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1666464484
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1666464484
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666464484
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1666464484
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1666464484
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1666464484
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1666464484
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1666464484
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1666464484
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1666464484
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1666464484
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1666464484
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1666464484
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1666464484
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1666464484
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1666464484
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1666464484
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1666464484
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1666464484
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1666464484
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1666464484
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1666464484
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1666464484
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1666464484
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1666464484
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1666464484
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1666464484
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1666464484
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1666464484
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1666464484
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1666464484
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1666464484
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666464484
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1666464484
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1666464484
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1666464484
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1666464484
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1666464484
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1666464484
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1666464484
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1666464484
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1666464484
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1666464484
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1666464484
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1666464484
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1666464484
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1666464484
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666464484
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666464484
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666464484
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666464484
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666464484
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666464484
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666464484
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666464484
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666464484
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666464484
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666464484
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666464484
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666464484
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666464484
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666464484
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666464484
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666464484
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1666464484
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1666464484
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1666464484
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1666464484
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1666464484
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1666464484
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1666464484
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1666464484
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1666464484
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1666464484
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1666464484
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1666464484
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1666464484
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1666464484
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1666464484
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1666464484
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1666464484
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1666464484
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1666464484
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1666464484
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1666464484
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1666464484
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1666464484
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1666464484
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1666464484
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1666464484
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1666464484
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1666464484
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1666464484
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1666464484
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1666464484
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1666464484
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666464484
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666464484
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666464484
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1666464484
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1666464484
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1666464484
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1666464484
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1666464484
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1666464484
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1666464484
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1666464484
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1666464484
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1666464484
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1666464484
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1666464484
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1666464484
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1666464484
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1666464484
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1666464484
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666464484
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666464484
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666464484
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666464484
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666464484
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666464484
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666464484
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666464484
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666464484
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666464484
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666464484
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666464484
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1666464484
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1666464484
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1666464484
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1666464484
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1666464484
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1666464484
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1666464484
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1666464484
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1666464484
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1666464484
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1666464484
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1666464484
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1666464484
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1666464484
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1666464484
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1666464484
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1666464484
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1666464484
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1666464484
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1666464484
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1666464484
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1666464484
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1666464484
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1666464484
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1666464484
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1666464484
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1666464484
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1666464484
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1666464484
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1666464484
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1666464484
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1666464484
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1666464484
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1666464484
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1666464484
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1666464484
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1666464484
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1666464484
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1666464484
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1666464484
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1666464484
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1666464484
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1666464484
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1666464484
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1666464484
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1666464484
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1666464484
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1666464484
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1666464484
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1666464484
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666464484
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666464484
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1666464484
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1666464484
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666464484
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1666464484
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666464484
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666464484
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666464484
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666464484
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666464484
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666464484
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666464484
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666464484
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666464484
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1666464484
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1666464484
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1666464484
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1666464484
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1666464484
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1666464484
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1666464484
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1666464484
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1666464484
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1666464484
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1666464484
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1666464484
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1666464484
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1666464484
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1666464484
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1666464484
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1666464484
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1666464484
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1666464484
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1666464484
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1666464484
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1666464484
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1666464484
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1666464484
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1666464484
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1666464484
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1666464484
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1666464484
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1666464484
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1666464484
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1666464484
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1666464484
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1666464484
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1666464484
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1666464484
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1666464484
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1666464484
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1666464484
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1666464484
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1666464484
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1666464484
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1666464484
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1666464484
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1666464484
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1666464484
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1666464484
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1666464484
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1666464484
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666464484
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1666464484
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666464484
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1666464484
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1666464484
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1666464484
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1666464484
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1666464484
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1666464484
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666464484
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666464484
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1666464484
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1666464484
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1666464484
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666464484
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1666464484
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1666464484
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1666464484
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1666464484
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1666464484
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1666464484
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1666464484
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1666464484
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1666464484
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1666464484
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1666464484
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1666464484
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1666464484
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1666464484
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1666464484
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1666464484
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1666464484
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1666464484
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1666464484
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1666464484
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1666464484
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1666464484
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1666464484
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666464484
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1666464484
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1666464484
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1666464484
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1666464484
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1666464484
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666464484
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1666464484
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1666464484
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1666464484
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1666464484
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1666464484
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1666464484
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1666464484
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1666464484
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1666464484
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1666464484
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1666464484
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1666464484
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1666464484
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1666464484
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1666464484
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1666464484
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1666464484
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1666464484
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1666464484
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_9
timestamp 1666464484
transform 1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1666464484
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666464484
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1666464484
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1666464484
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1666464484
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1666464484
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1666464484
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1666464484
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1666464484
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1666464484
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1666464484
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1666464484
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1666464484
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1666464484
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1666464484
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1666464484
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1666464484
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1666464484
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1666464484
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1666464484
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1666464484
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1666464484
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1666464484
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1666464484
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1666464484
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1666464484
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1666464484
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1666464484
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1666464484
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1666464484
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1666464484
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1666464484
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1666464484
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1666464484
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1666464484
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1666464484
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1666464484
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666464484
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1666464484
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1666464484
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1666464484
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1666464484
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1666464484
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1666464484
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1666464484
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1666464484
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1666464484
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1666464484
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1666464484
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1666464484
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1666464484
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1666464484
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1666464484
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1666464484
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1666464484
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1666464484
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1666464484
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1666464484
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1666464484
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1666464484
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1666464484
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1666464484
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1666464484
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1666464484
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1666464484
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1666464484
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1666464484
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1666464484
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1666464484
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1666464484
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1666464484
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1666464484
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1666464484
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1666464484
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1666464484
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1666464484
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1666464484
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1666464484
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1666464484
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1666464484
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1666464484
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1666464484
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1666464484
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1666464484
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1666464484
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1666464484
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1666464484
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1666464484
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1666464484
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1666464484
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1666464484
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1666464484
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1666464484
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1666464484
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1666464484
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1666464484
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1666464484
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1666464484
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1666464484
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1666464484
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1666464484
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1666464484
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1666464484
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1666464484
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1666464484
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1666464484
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1666464484
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1666464484
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1666464484
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1666464484
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1666464484
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1666464484
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1666464484
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1666464484
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1666464484
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1666464484
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1666464484
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1666464484
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1666464484
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1666464484
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1666464484
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1666464484
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1666464484
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1666464484
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1666464484
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1666464484
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1666464484
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1666464484
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1666464484
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1666464484
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1666464484
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1666464484
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1666464484
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1666464484
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1666464484
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1666464484
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1666464484
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1666464484
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1666464484
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1666464484
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1666464484
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1666464484
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1666464484
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1666464484
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1666464484
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1666464484
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1666464484
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1666464484
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1666464484
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1666464484
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1666464484
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1666464484
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1666464484
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1666464484
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1666464484
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1666464484
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1666464484
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1666464484
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1666464484
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1666464484
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1666464484
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1666464484
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1666464484
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1666464484
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1666464484
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1666464484
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1666464484
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1666464484
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1666464484
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1666464484
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1666464484
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1666464484
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1666464484
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1666464484
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1666464484
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1666464484
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1666464484
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1666464484
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1666464484
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1666464484
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1666464484
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1666464484
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1666464484
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1666464484
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1666464484
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1666464484
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1666464484
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1666464484
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1666464484
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1666464484
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1666464484
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1666464484
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1666464484
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1666464484
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1666464484
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1666464484
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1666464484
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1666464484
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1666464484
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1666464484
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1666464484
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1666464484
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1666464484
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1666464484
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1666464484
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1666464484
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1666464484
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1666464484
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1666464484
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1666464484
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1666464484
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1666464484
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1666464484
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1666464484
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1666464484
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1666464484
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1666464484
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1666464484
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1666464484
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1666464484
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1666464484
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1666464484
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1666464484
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1666464484
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1666464484
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1666464484
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1666464484
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1666464484
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1666464484
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1666464484
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1666464484
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1666464484
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1666464484
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1666464484
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1666464484
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1666464484
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1666464484
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1666464484
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1666464484
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1666464484
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1666464484
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1666464484
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1666464484
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1666464484
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1666464484
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1666464484
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1666464484
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1666464484
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1666464484
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1666464484
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1666464484
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1666464484
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1666464484
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1666464484
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1666464484
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1666464484
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1666464484
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_609
timestamp 1666464484
transform 1 0 57132 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_614
timestamp 1666464484
transform 1 0 57592 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_617
timestamp 1666464484
transform 1 0 57868 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_623
timestamp 1666464484
transform 1 0 58420 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1666464484
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1666464484
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1666464484
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1666464484
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1666464484
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1666464484
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1666464484
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1666464484
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1666464484
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1666464484
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1666464484
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1666464484
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1666464484
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1666464484
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1666464484
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1666464484
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1666464484
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1666464484
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1666464484
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1666464484
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1666464484
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1666464484
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1666464484
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1666464484
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1666464484
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1666464484
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1666464484
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1666464484
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1666464484
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1666464484
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1666464484
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1666464484
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1666464484
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1666464484
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1666464484
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1666464484
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1666464484
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1666464484
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1666464484
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1666464484
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1666464484
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1666464484
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1666464484
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1666464484
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1666464484
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1666464484
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1666464484
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1666464484
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1666464484
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1666464484
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1666464484
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1666464484
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1666464484
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1666464484
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1666464484
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1666464484
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1666464484
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1666464484
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1666464484
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1666464484
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1666464484
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1666464484
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1666464484
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1666464484
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1666464484
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1666464484
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1666464484
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1666464484
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1666464484
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1666464484
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1666464484
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1666464484
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1666464484
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1666464484
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1666464484
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1666464484
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1666464484
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1666464484
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1666464484
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1666464484
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1666464484
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1666464484
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1666464484
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1666464484
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1666464484
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1666464484
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1666464484
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1666464484
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1666464484
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1666464484
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1666464484
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1666464484
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1666464484
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1666464484
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1666464484
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1666464484
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1666464484
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1666464484
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1666464484
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1666464484
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1666464484
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1666464484
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1666464484
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1666464484
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1666464484
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1666464484
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1666464484
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1666464484
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1666464484
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1666464484
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1666464484
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1666464484
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1666464484
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1666464484
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1666464484
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1666464484
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1666464484
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1666464484
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1666464484
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1666464484
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1666464484
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1666464484
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1666464484
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1666464484
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1666464484
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1666464484
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1666464484
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1666464484
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1666464484
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1666464484
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1666464484
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1666464484
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1666464484
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1666464484
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1666464484
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1666464484
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1666464484
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1666464484
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1666464484
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1666464484
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1666464484
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1666464484
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1666464484
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1666464484
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1666464484
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1666464484
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1666464484
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1666464484
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1666464484
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1666464484
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1666464484
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1666464484
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1666464484
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1666464484
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1666464484
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1666464484
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1666464484
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1666464484
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1666464484
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1666464484
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1666464484
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1666464484
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1666464484
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1666464484
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1666464484
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1666464484
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1666464484
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1666464484
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1666464484
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1666464484
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1666464484
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1666464484
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1666464484
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1666464484
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1666464484
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1666464484
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1666464484
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1666464484
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1666464484
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1666464484
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1666464484
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1666464484
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1666464484
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1666464484
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1666464484
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1666464484
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1666464484
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1666464484
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1666464484
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1666464484
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1666464484
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1666464484
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1666464484
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1666464484
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1666464484
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1666464484
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1666464484
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1666464484
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1666464484
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1666464484
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1666464484
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1666464484
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1666464484
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1666464484
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1666464484
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1666464484
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1666464484
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1666464484
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1666464484
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1666464484
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1666464484
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1666464484
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1666464484
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1666464484
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1666464484
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1666464484
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1666464484
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1666464484
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1666464484
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1666464484
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1666464484
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1666464484
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1666464484
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1666464484
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1666464484
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1666464484
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1666464484
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1666464484
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1666464484
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1666464484
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1666464484
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1666464484
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1666464484
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1666464484
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1666464484
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1666464484
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1666464484
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1666464484
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1666464484
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1666464484
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1666464484
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1666464484
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1666464484
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1666464484
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1666464484
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1666464484
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1666464484
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1666464484
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1666464484
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1666464484
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1666464484
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1666464484
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1666464484
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1666464484
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1666464484
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1666464484
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1666464484
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1666464484
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1666464484
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1666464484
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1666464484
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1666464484
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1666464484
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1666464484
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1666464484
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1666464484
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1666464484
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1666464484
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1666464484
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1666464484
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1666464484
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1666464484
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1666464484
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1666464484
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1666464484
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1666464484
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1666464484
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1666464484
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1666464484
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1666464484
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1666464484
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1666464484
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1666464484
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1666464484
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1666464484
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1666464484
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1666464484
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1666464484
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1666464484
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1666464484
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1666464484
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1666464484
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1666464484
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1666464484
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1666464484
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1666464484
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1666464484
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1666464484
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1666464484
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1666464484
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1666464484
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1666464484
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1666464484
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1666464484
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1666464484
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1666464484
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1666464484
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1666464484
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1666464484
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1666464484
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1666464484
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1666464484
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1666464484
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1666464484
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1666464484
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1666464484
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1666464484
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1666464484
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1666464484
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1666464484
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1666464484
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1666464484
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1666464484
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1666464484
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1666464484
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1666464484
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1666464484
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1666464484
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1666464484
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1666464484
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1666464484
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1666464484
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1666464484
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1666464484
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1666464484
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1666464484
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1666464484
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1666464484
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1666464484
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1666464484
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1666464484
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1666464484
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1666464484
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1666464484
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1666464484
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1666464484
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1666464484
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1666464484
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1666464484
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1666464484
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1666464484
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1666464484
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1666464484
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1666464484
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1666464484
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1666464484
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1666464484
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1666464484
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1666464484
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1666464484
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1666464484
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1666464484
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1666464484
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1666464484
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1666464484
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1666464484
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1666464484
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1666464484
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1666464484
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1666464484
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1666464484
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1666464484
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1666464484
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1666464484
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1666464484
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1666464484
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1666464484
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1666464484
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1666464484
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1666464484
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1666464484
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1666464484
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1666464484
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1666464484
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1666464484
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1666464484
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1666464484
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1666464484
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1666464484
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1666464484
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1666464484
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1666464484
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1666464484
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1666464484
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1666464484
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1666464484
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1666464484
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1666464484
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1666464484
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1666464484
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1666464484
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1666464484
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1666464484
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1666464484
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1666464484
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1666464484
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1666464484
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1666464484
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1666464484
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1666464484
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1666464484
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1666464484
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1666464484
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1666464484
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1666464484
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1666464484
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1666464484
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1666464484
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1666464484
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1666464484
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1666464484
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1666464484
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1666464484
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1666464484
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1666464484
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1666464484
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1666464484
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1666464484
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1666464484
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1666464484
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1666464484
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1666464484
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1666464484
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1666464484
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1666464484
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1666464484
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1666464484
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1666464484
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1666464484
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1666464484
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1666464484
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1666464484
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1666464484
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1666464484
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1666464484
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1666464484
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1666464484
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1666464484
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1666464484
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1666464484
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1666464484
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1666464484
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1666464484
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1666464484
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1666464484
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1666464484
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1666464484
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1666464484
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1666464484
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1666464484
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1666464484
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1666464484
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1666464484
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1666464484
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1666464484
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1666464484
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1666464484
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1666464484
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1666464484
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1666464484
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1666464484
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1666464484
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1666464484
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1666464484
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1666464484
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1666464484
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1666464484
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1666464484
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1666464484
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1666464484
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1666464484
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1666464484
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1666464484
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1666464484
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1666464484
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1666464484
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1666464484
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1666464484
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1666464484
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1666464484
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1666464484
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1666464484
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1666464484
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1666464484
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1666464484
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1666464484
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1666464484
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1666464484
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1666464484
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1666464484
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1666464484
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1666464484
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1666464484
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1666464484
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1666464484
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1666464484
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1666464484
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1666464484
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1666464484
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1666464484
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1666464484
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1666464484
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_9
timestamp 1666464484
transform 1 0 1932 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1666464484
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1666464484
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1666464484
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1666464484
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1666464484
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1666464484
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1666464484
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1666464484
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1666464484
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1666464484
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1666464484
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1666464484
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1666464484
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1666464484
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1666464484
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1666464484
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1666464484
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1666464484
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1666464484
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1666464484
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1666464484
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1666464484
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1666464484
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1666464484
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1666464484
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1666464484
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1666464484
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1666464484
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1666464484
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1666464484
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1666464484
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1666464484
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1666464484
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1666464484
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1666464484
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1666464484
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1666464484
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1666464484
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1666464484
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1666464484
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1666464484
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1666464484
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1666464484
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1666464484
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1666464484
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1666464484
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1666464484
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1666464484
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1666464484
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1666464484
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1666464484
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1666464484
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1666464484
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1666464484
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1666464484
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1666464484
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1666464484
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1666464484
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1666464484
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1666464484
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1666464484
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1666464484
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1666464484
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1666464484
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1666464484
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1666464484
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1666464484
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1666464484
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1666464484
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1666464484
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1666464484
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1666464484
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1666464484
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1666464484
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1666464484
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1666464484
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1666464484
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1666464484
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1666464484
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1666464484
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1666464484
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1666464484
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1666464484
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1666464484
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1666464484
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1666464484
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1666464484
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1666464484
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1666464484
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1666464484
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1666464484
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1666464484
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1666464484
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1666464484
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1666464484
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1666464484
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1666464484
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1666464484
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1666464484
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1666464484
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1666464484
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1666464484
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1666464484
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1666464484
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1666464484
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1666464484
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1666464484
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1666464484
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1666464484
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1666464484
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1666464484
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1666464484
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1666464484
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1666464484
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1666464484
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1666464484
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1666464484
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1666464484
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1666464484
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1666464484
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1666464484
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1666464484
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1666464484
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1666464484
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1666464484
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1666464484
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1666464484
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1666464484
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1666464484
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1666464484
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1666464484
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1666464484
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1666464484
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1666464484
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1666464484
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1666464484
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1666464484
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1666464484
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1666464484
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1666464484
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1666464484
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1666464484
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1666464484
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1666464484
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1666464484
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1666464484
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1666464484
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1666464484
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1666464484
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1666464484
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1666464484
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1666464484
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1666464484
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1666464484
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1666464484
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1666464484
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1666464484
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1666464484
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1666464484
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1666464484
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1666464484
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1666464484
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1666464484
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1666464484
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1666464484
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1666464484
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1666464484
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1666464484
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1666464484
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1666464484
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1666464484
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1666464484
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1666464484
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1666464484
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1666464484
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1666464484
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1666464484
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1666464484
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1666464484
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1666464484
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1666464484
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1666464484
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1666464484
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1666464484
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1666464484
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1666464484
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1666464484
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1666464484
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1666464484
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1666464484
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1666464484
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1666464484
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1666464484
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1666464484
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1666464484
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_615
timestamp 1666464484
transform 1 0 57684 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_623
timestamp 1666464484
transform 1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1666464484
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1666464484
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1666464484
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1666464484
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1666464484
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1666464484
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1666464484
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1666464484
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1666464484
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1666464484
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1666464484
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1666464484
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1666464484
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1666464484
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1666464484
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1666464484
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1666464484
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1666464484
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1666464484
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1666464484
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1666464484
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1666464484
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1666464484
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1666464484
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1666464484
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1666464484
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1666464484
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1666464484
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1666464484
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1666464484
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1666464484
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1666464484
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1666464484
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1666464484
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1666464484
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1666464484
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1666464484
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1666464484
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1666464484
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1666464484
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1666464484
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1666464484
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1666464484
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1666464484
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1666464484
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1666464484
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1666464484
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1666464484
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1666464484
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1666464484
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1666464484
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1666464484
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1666464484
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1666464484
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1666464484
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1666464484
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1666464484
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1666464484
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1666464484
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1666464484
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1666464484
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1666464484
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1666464484
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1666464484
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1666464484
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1666464484
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1666464484
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1666464484
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1666464484
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1666464484
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1666464484
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1666464484
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1666464484
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1666464484
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1666464484
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1666464484
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1666464484
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1666464484
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1666464484
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1666464484
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1666464484
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1666464484
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1666464484
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1666464484
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1666464484
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1666464484
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1666464484
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1666464484
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1666464484
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1666464484
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1666464484
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1666464484
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1666464484
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1666464484
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1666464484
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1666464484
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1666464484
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1666464484
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1666464484
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1666464484
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1666464484
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1666464484
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1666464484
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1666464484
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1666464484
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1666464484
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1666464484
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1666464484
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1666464484
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1666464484
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1666464484
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1666464484
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1666464484
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1666464484
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1666464484
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1666464484
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1666464484
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1666464484
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1666464484
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1666464484
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1666464484
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1666464484
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1666464484
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1666464484
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1666464484
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1666464484
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1666464484
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1666464484
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1666464484
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1666464484
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1666464484
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1666464484
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1666464484
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1666464484
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1666464484
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1666464484
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1666464484
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1666464484
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1666464484
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1666464484
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1666464484
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1666464484
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1666464484
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1666464484
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1666464484
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1666464484
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1666464484
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1666464484
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1666464484
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1666464484
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1666464484
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1666464484
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1666464484
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1666464484
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1666464484
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1666464484
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1666464484
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1666464484
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1666464484
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1666464484
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1666464484
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1666464484
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1666464484
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1666464484
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1666464484
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1666464484
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1666464484
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1666464484
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1666464484
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1666464484
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1666464484
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1666464484
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1666464484
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1666464484
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1666464484
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1666464484
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1666464484
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1666464484
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1666464484
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1666464484
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1666464484
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1666464484
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1666464484
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1666464484
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1666464484
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1666464484
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1666464484
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1666464484
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1666464484
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1666464484
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1666464484
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1666464484
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1666464484
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1666464484
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1666464484
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_617
timestamp 1666464484
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1666464484
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1666464484
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1666464484
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1666464484
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1666464484
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1666464484
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1666464484
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1666464484
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1666464484
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1666464484
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1666464484
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1666464484
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1666464484
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1666464484
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1666464484
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_153
timestamp 1666464484
transform 1 0 15180 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_163
timestamp 1666464484
transform 1 0 16100 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_175
timestamp 1666464484
transform 1 0 17204 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_187
timestamp 1666464484
transform 1 0 18308 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1666464484
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1666464484
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1666464484
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1666464484
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1666464484
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1666464484
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1666464484
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1666464484
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1666464484
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1666464484
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1666464484
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1666464484
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1666464484
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1666464484
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1666464484
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1666464484
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1666464484
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1666464484
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1666464484
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1666464484
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1666464484
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1666464484
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1666464484
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1666464484
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1666464484
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1666464484
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_433
timestamp 1666464484
transform 1 0 40940 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_438
timestamp 1666464484
transform 1 0 41400 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_444
timestamp 1666464484
transform 1 0 41952 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_456
timestamp 1666464484
transform 1 0 43056 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_468
timestamp 1666464484
transform 1 0 44160 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1666464484
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1666464484
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1666464484
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1666464484
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_527
timestamp 1666464484
transform 1 0 49588 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1666464484
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1666464484
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1666464484
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1666464484
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1666464484
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1666464484
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1666464484
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1666464484
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1666464484
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1666464484
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_9
timestamp 1666464484
transform 1 0 1932 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1666464484
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1666464484
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_29
timestamp 1666464484
transform 1 0 3772 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_35
timestamp 1666464484
transform 1 0 4324 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_41
timestamp 1666464484
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1666464484
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1666464484
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1666464484
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_81
timestamp 1666464484
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_85
timestamp 1666464484
transform 1 0 8924 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_93
timestamp 1666464484
transform 1 0 9660 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_98
timestamp 1666464484
transform 1 0 10120 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_104
timestamp 1666464484
transform 1 0 10672 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1666464484
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1666464484
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_137
timestamp 1666464484
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_141
timestamp 1666464484
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_153
timestamp 1666464484
transform 1 0 15180 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1666464484
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1666464484
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1666464484
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1666464484
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1666464484
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_197
timestamp 1666464484
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_209
timestamp 1666464484
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_221
timestamp 1666464484
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_225
timestamp 1666464484
transform 1 0 21804 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_231
timestamp 1666464484
transform 1 0 22356 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1666464484
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_249
timestamp 1666464484
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_253
timestamp 1666464484
transform 1 0 24380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_265
timestamp 1666464484
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_277
timestamp 1666464484
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_281
timestamp 1666464484
transform 1 0 26956 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_287
timestamp 1666464484
transform 1 0 27508 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1666464484
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_305
timestamp 1666464484
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_309
timestamp 1666464484
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_321
timestamp 1666464484
transform 1 0 30636 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_329
timestamp 1666464484
transform 1 0 31372 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_334
timestamp 1666464484
transform 1 0 31832 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_337
timestamp 1666464484
transform 1 0 32108 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_345
timestamp 1666464484
transform 1 0 32844 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_357
timestamp 1666464484
transform 1 0 33948 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_363
timestamp 1666464484
transform 1 0 34500 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_365
timestamp 1666464484
transform 1 0 34684 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_377
timestamp 1666464484
transform 1 0 35788 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_389
timestamp 1666464484
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_101_393
timestamp 1666464484
transform 1 0 37260 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_398
timestamp 1666464484
transform 1 0 37720 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_406
timestamp 1666464484
transform 1 0 38456 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_418
timestamp 1666464484
transform 1 0 39560 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_421
timestamp 1666464484
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_433
timestamp 1666464484
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1666464484
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_449
timestamp 1666464484
transform 1 0 42412 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_457
timestamp 1666464484
transform 1 0 43148 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_462
timestamp 1666464484
transform 1 0 43608 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_468
timestamp 1666464484
transform 1 0 44160 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_477
timestamp 1666464484
transform 1 0 44988 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_489
timestamp 1666464484
transform 1 0 46092 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_501
timestamp 1666464484
transform 1 0 47196 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1666464484
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_517
timestamp 1666464484
transform 1 0 48668 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_525
timestamp 1666464484
transform 1 0 49404 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_531
timestamp 1666464484
transform 1 0 49956 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_533
timestamp 1666464484
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_545
timestamp 1666464484
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_557
timestamp 1666464484
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1666464484
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1666464484
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1666464484
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_589
timestamp 1666464484
transform 1 0 55292 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_595
timestamp 1666464484
transform 1 0 55844 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_607
timestamp 1666464484
transform 1 0 56948 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_611
timestamp 1666464484
transform 1 0 57316 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_614
timestamp 1666464484
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_617
timestamp 1666464484
transform 1 0 57868 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_623
timestamp 1666464484
transform 1 0 58420 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0985_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 53544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0986_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 52440 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0987_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 54464 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0988_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 54188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0989_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 54004 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1666464484
transform -1 0 56488 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0991_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 55844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0992_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 52440 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _0993_
timestamp 1666464484
transform -1 0 55016 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0994_
timestamp 1666464484
transform -1 0 53452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_4  _0995_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 55476 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _0996_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 52348 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0997_
timestamp 1666464484
transform 1 0 54096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_2  _0998_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 56212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_4  _0999_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 57132 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__a2111oi_4  _1000_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 55200 0 -1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_4  _1001_
timestamp 1666464484
transform 1 0 39008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1002_
timestamp 1666464484
transform -1 0 39928 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1003_
timestamp 1666464484
transform -1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1004_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 42964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _1005_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1006_
timestamp 1666464484
transform 1 0 35052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1007_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1008_
timestamp 1666464484
transform -1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_2  _1009_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1010_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 40480 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1011_
timestamp 1666464484
transform 1 0 41400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1012_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37628 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1013_
timestamp 1666464484
transform -1 0 31832 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1014_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 39376 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1015_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1016_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1017_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 32936 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _1018_
timestamp 1666464484
transform 1 0 26680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1019_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1020_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31832 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1666464484
transform -1 0 22632 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1022_
timestamp 1666464484
transform -1 0 44068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1023_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43240 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1024_
timestamp 1666464484
transform 1 0 42780 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1025_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 42872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1666464484
transform 1 0 24564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1027_
timestamp 1666464484
transform 1 0 24564 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1666464484
transform 1 0 23644 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1666464484
transform 1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1030_
timestamp 1666464484
transform 1 0 41952 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1666464484
transform -1 0 42872 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1032_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 22724 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1666464484
transform -1 0 22632 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1034_
timestamp 1666464484
transform 1 0 26404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1035_
timestamp 1666464484
transform 1 0 32292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1666464484
transform 1 0 24288 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1037_
timestamp 1666464484
transform 1 0 24748 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1038_
timestamp 1666464484
transform 1 0 29992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1039_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33580 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1040_
timestamp 1666464484
transform 1 0 30084 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1041_
timestamp 1666464484
transform -1 0 35328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1042_
timestamp 1666464484
transform 1 0 37444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1043_
timestamp 1666464484
transform -1 0 29256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1044_
timestamp 1666464484
transform -1 0 31280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1666464484
transform 1 0 29716 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1046_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28704 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1047_
timestamp 1666464484
transform 1 0 30820 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1048_
timestamp 1666464484
transform -1 0 26588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_2  _1049_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33304 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_2  _1050_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1051_
timestamp 1666464484
transform 1 0 29716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30176 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1053_
timestamp 1666464484
transform -1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1054_
timestamp 1666464484
transform -1 0 39284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1055_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1666464484
transform 1 0 36708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1057_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 41952 0 -1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_1  _1058_
timestamp 1666464484
transform 1 0 30176 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_2  _1059_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30360 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1060_
timestamp 1666464484
transform 1 0 27508 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1061_
timestamp 1666464484
transform 1 0 28704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _1062_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1063_
timestamp 1666464484
transform -1 0 25024 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1666464484
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1065_
timestamp 1666464484
transform -1 0 38364 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1066_
timestamp 1666464484
transform 1 0 28612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1067_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34408 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _1068_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26680 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 1666464484
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1070_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27600 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1071_
timestamp 1666464484
transform 1 0 25392 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1072_
timestamp 1666464484
transform -1 0 31096 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1073_
timestamp 1666464484
transform 1 0 24932 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1074_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1075_
timestamp 1666464484
transform -1 0 29900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1076_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1077_
timestamp 1666464484
transform 1 0 25668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1078_
timestamp 1666464484
transform 1 0 26220 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1666464484
transform -1 0 35788 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1080_
timestamp 1666464484
transform -1 0 35512 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1081_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_2  _1082_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1666464484
transform 1 0 31924 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1084_
timestamp 1666464484
transform 1 0 38272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _1085_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 32936 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1086_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 38272 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1087_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1088_
timestamp 1666464484
transform 1 0 24748 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2b_4  _1089_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35972 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__a21oi_1  _1090_
timestamp 1666464484
transform -1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1091_
timestamp 1666464484
transform 1 0 30820 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1092_
timestamp 1666464484
transform -1 0 31188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1093_
timestamp 1666464484
transform -1 0 33120 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _1094_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _1095_
timestamp 1666464484
transform 1 0 27140 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1096_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25484 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1097_
timestamp 1666464484
transform 1 0 27508 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1098_
timestamp 1666464484
transform 1 0 27692 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1666464484
transform -1 0 25668 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1100_
timestamp 1666464484
transform 1 0 25484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1101_
timestamp 1666464484
transform 1 0 25392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1102_
timestamp 1666464484
transform 1 0 25116 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _1103_
timestamp 1666464484
transform 1 0 31188 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _1104_
timestamp 1666464484
transform 1 0 25760 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1105_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 38732 0 1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1666464484
transform -1 0 25668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1107_
timestamp 1666464484
transform 1 0 35144 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1108_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34408 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1109_
timestamp 1666464484
transform 1 0 27968 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1110_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1111_
timestamp 1666464484
transform -1 0 27876 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1112_
timestamp 1666464484
transform -1 0 26312 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1113_
timestamp 1666464484
transform 1 0 25392 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1114_
timestamp 1666464484
transform -1 0 31556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1115_
timestamp 1666464484
transform -1 0 28888 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1116_
timestamp 1666464484
transform -1 0 27508 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1117_
timestamp 1666464484
transform -1 0 27692 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _1118_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32384 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_1  _1119_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1120_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34408 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1121_
timestamp 1666464484
transform 1 0 28244 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1122_
timestamp 1666464484
transform 1 0 27784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1123_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1124_
timestamp 1666464484
transform -1 0 27876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1125_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26220 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1126_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_2  _1127_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30268 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1128_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29900 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__o31a_1  _1129_
timestamp 1666464484
transform 1 0 28704 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1130_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37996 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1131_
timestamp 1666464484
transform -1 0 40388 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1132_
timestamp 1666464484
transform 1 0 28428 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1133_
timestamp 1666464484
transform -1 0 29992 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1134_
timestamp 1666464484
transform -1 0 28336 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _1135_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27324 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1136_
timestamp 1666464484
transform 1 0 27140 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1137_
timestamp 1666464484
transform 1 0 26220 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1138_
timestamp 1666464484
transform -1 0 26680 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1139_
timestamp 1666464484
transform -1 0 27692 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_2  _1140_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25300 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1141_
timestamp 1666464484
transform 1 0 24564 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 1666464484
transform -1 0 30360 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _1143_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1144_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1145_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28060 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1146_
timestamp 1666464484
transform -1 0 25024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1147_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25024 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1148_
timestamp 1666464484
transform 1 0 25392 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1149_
timestamp 1666464484
transform -1 0 29532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1150_
timestamp 1666464484
transform 1 0 28796 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _1151_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1152_
timestamp 1666464484
transform -1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1153_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25944 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1154_
timestamp 1666464484
transform 1 0 26036 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1155_
timestamp 1666464484
transform -1 0 24104 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _1156_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26680 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1666464484
transform 1 0 30452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1158_
timestamp 1666464484
transform -1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1159_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26496 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _1160_
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1161_
timestamp 1666464484
transform 1 0 31464 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1162_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25668 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _1163_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24932 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1164_
timestamp 1666464484
transform 1 0 28704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1165_
timestamp 1666464484
transform -1 0 30176 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1166_
timestamp 1666464484
transform -1 0 32936 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1167_
timestamp 1666464484
transform 1 0 29716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1168_
timestamp 1666464484
transform 1 0 29716 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1169_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31464 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1170_
timestamp 1666464484
transform -1 0 31096 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1171_
timestamp 1666464484
transform 1 0 30268 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1172_
timestamp 1666464484
transform -1 0 29256 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1173_
timestamp 1666464484
transform -1 0 29256 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1174_
timestamp 1666464484
transform 1 0 28704 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1175_
timestamp 1666464484
transform -1 0 29716 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1176_
timestamp 1666464484
transform -1 0 26404 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1177_
timestamp 1666464484
transform 1 0 25944 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1178_
timestamp 1666464484
transform 1 0 23736 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1179_
timestamp 1666464484
transform 1 0 24564 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1180_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24380 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1181_
timestamp 1666464484
transform 1 0 24564 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1182_
timestamp 1666464484
transform -1 0 25668 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1183_
timestamp 1666464484
transform -1 0 25760 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_1  _1184_
timestamp 1666464484
transform -1 0 25116 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1185_
timestamp 1666464484
transform 1 0 24288 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1186_
timestamp 1666464484
transform 1 0 23736 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1187_
timestamp 1666464484
transform -1 0 25024 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1188_
timestamp 1666464484
transform -1 0 24104 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1189_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 24104 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1190_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 23736 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__o32ai_4  _1191_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26036 0 1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__and2b_1  _1192_
timestamp 1666464484
transform -1 0 23644 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1193_
timestamp 1666464484
transform -1 0 23644 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_1  _1194_
timestamp 1666464484
transform 1 0 26496 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1195_
timestamp 1666464484
transform 1 0 26036 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1196_
timestamp 1666464484
transform 1 0 26128 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1197_
timestamp 1666464484
transform -1 0 29992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1198_
timestamp 1666464484
transform 1 0 28244 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1199_
timestamp 1666464484
transform 1 0 28244 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1200_
timestamp 1666464484
transform -1 0 33948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1201_
timestamp 1666464484
transform 1 0 33764 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1202_
timestamp 1666464484
transform 1 0 35604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1203_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34224 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1204_
timestamp 1666464484
transform 1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1205_
timestamp 1666464484
transform 1 0 25300 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1206_
timestamp 1666464484
transform 1 0 24564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1207_
timestamp 1666464484
transform -1 0 25024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1208_
timestamp 1666464484
transform -1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1209_
timestamp 1666464484
transform 1 0 27232 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1210_
timestamp 1666464484
transform -1 0 29256 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1211_
timestamp 1666464484
transform -1 0 26680 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1212_
timestamp 1666464484
transform 1 0 27784 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1213_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1214_
timestamp 1666464484
transform 1 0 27140 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1215_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1216_
timestamp 1666464484
transform -1 0 28060 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1217_
timestamp 1666464484
transform 1 0 27324 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1218_
timestamp 1666464484
transform -1 0 28428 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1219_
timestamp 1666464484
transform 1 0 27968 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1220_
timestamp 1666464484
transform 1 0 27600 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1221_
timestamp 1666464484
transform 1 0 28060 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1222_
timestamp 1666464484
transform -1 0 32568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1223_
timestamp 1666464484
transform -1 0 30912 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1224_
timestamp 1666464484
transform 1 0 29440 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1225_
timestamp 1666464484
transform -1 0 29992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1226_
timestamp 1666464484
transform -1 0 30176 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1227_
timestamp 1666464484
transform -1 0 29256 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_1  _1228_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29348 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 1666464484
transform 1 0 29992 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1230_
timestamp 1666464484
transform -1 0 28336 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1231_
timestamp 1666464484
transform -1 0 28336 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1232_
timestamp 1666464484
transform -1 0 27600 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _1233_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27968 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1234_
timestamp 1666464484
transform -1 0 28980 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1235_
timestamp 1666464484
transform 1 0 24472 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _1236_
timestamp 1666464484
transform -1 0 25208 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1237_
timestamp 1666464484
transform -1 0 25760 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1238_
timestamp 1666464484
transform 1 0 31556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 1666464484
transform -1 0 32660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1240_
timestamp 1666464484
transform -1 0 33304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1241_
timestamp 1666464484
transform -1 0 34224 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1242_
timestamp 1666464484
transform 1 0 34868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1243_
timestamp 1666464484
transform -1 0 33396 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1244_
timestamp 1666464484
transform 1 0 33580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1245_
timestamp 1666464484
transform 1 0 33764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1246_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32752 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1247_
timestamp 1666464484
transform -1 0 31740 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 1666464484
transform -1 0 31832 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1249_
timestamp 1666464484
transform -1 0 32016 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1250_
timestamp 1666464484
transform -1 0 26588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1251_
timestamp 1666464484
transform 1 0 31004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1252_
timestamp 1666464484
transform -1 0 31372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1253_
timestamp 1666464484
transform -1 0 31832 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1254_
timestamp 1666464484
transform 1 0 31372 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1255_
timestamp 1666464484
transform -1 0 30636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1256_
timestamp 1666464484
transform -1 0 31740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1257_
timestamp 1666464484
transform -1 0 31464 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1258_
timestamp 1666464484
transform 1 0 30728 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1259_
timestamp 1666464484
transform 1 0 30544 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _1260_
timestamp 1666464484
transform 1 0 29716 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1261_
timestamp 1666464484
transform -1 0 31280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1262_
timestamp 1666464484
transform 1 0 30728 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _1263_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31832 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1264_
timestamp 1666464484
transform -1 0 32936 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1265_
timestamp 1666464484
transform 1 0 33488 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1266_
timestamp 1666464484
transform 1 0 32476 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1267_
timestamp 1666464484
transform -1 0 38272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 1666464484
transform -1 0 38272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1269_
timestamp 1666464484
transform 1 0 30360 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1270_
timestamp 1666464484
transform -1 0 31372 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1271_
timestamp 1666464484
transform 1 0 30728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1272_
timestamp 1666464484
transform 1 0 28980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1273_
timestamp 1666464484
transform -1 0 30084 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1274_
timestamp 1666464484
transform 1 0 30176 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1275_
timestamp 1666464484
transform 1 0 31188 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _1276_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31004 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1277_
timestamp 1666464484
transform 1 0 27876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1278_
timestamp 1666464484
transform 1 0 28428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1279_
timestamp 1666464484
transform 1 0 29808 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _1280_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30728 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o2111ai_4  _1281_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31372 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__o21a_1  _1282_
timestamp 1666464484
transform -1 0 29072 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1283_
timestamp 1666464484
transform 1 0 29716 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1284_
timestamp 1666464484
transform 1 0 29992 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1285_
timestamp 1666464484
transform 1 0 58144 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1666464484
transform 1 0 32200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1287_
timestamp 1666464484
transform 1 0 34500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1288_
timestamp 1666464484
transform 1 0 35328 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1289_
timestamp 1666464484
transform 1 0 32292 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1290_
timestamp 1666464484
transform 1 0 40020 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1291_
timestamp 1666464484
transform 1 0 32292 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1292_
timestamp 1666464484
transform 1 0 32016 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1293_
timestamp 1666464484
transform -1 0 33028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1294_
timestamp 1666464484
transform 1 0 32476 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1295_
timestamp 1666464484
transform 1 0 32384 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1296_
timestamp 1666464484
transform 1 0 33396 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1297_
timestamp 1666464484
transform 1 0 33672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1298_
timestamp 1666464484
transform 1 0 33396 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1299_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1300_
timestamp 1666464484
transform -1 0 33028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1301_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 33212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1302_
timestamp 1666464484
transform 1 0 32936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1303_
timestamp 1666464484
transform -1 0 33304 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _1304_
timestamp 1666464484
transform -1 0 31740 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1305_
timestamp 1666464484
transform 1 0 33672 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1306_
timestamp 1666464484
transform 1 0 33580 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1307_
timestamp 1666464484
transform -1 0 33856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1308_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 33672 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1309_
timestamp 1666464484
transform 1 0 32936 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_1  _1310_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29532 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1311_
timestamp 1666464484
transform -1 0 35696 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1312_
timestamp 1666464484
transform -1 0 39376 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1313_
timestamp 1666464484
transform 1 0 37444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1314_
timestamp 1666464484
transform 1 0 36524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1315_
timestamp 1666464484
transform -1 0 38916 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1316_
timestamp 1666464484
transform 1 0 35972 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a311oi_4  _1317_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35328 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1318_
timestamp 1666464484
transform -1 0 35696 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1319_
timestamp 1666464484
transform -1 0 33948 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1320_
timestamp 1666464484
transform 1 0 30728 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1321_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31832 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1322_
timestamp 1666464484
transform 1 0 30728 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1323_
timestamp 1666464484
transform 1 0 31372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1324_
timestamp 1666464484
transform 1 0 31280 0 1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1325_
timestamp 1666464484
transform 1 0 37904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _1326_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1327_
timestamp 1666464484
transform 1 0 39192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1328_
timestamp 1666464484
transform 1 0 39008 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1329_
timestamp 1666464484
transform -1 0 40296 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1330_
timestamp 1666464484
transform -1 0 37996 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1331_
timestamp 1666464484
transform 1 0 37536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1332_
timestamp 1666464484
transform 1 0 38088 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1333_
timestamp 1666464484
transform -1 0 40848 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1334_
timestamp 1666464484
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1335_
timestamp 1666464484
transform 1 0 39836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1336_
timestamp 1666464484
transform 1 0 40020 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1337_
timestamp 1666464484
transform -1 0 40572 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1338_
timestamp 1666464484
transform 1 0 39100 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1339_
timestamp 1666464484
transform 1 0 39560 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1340_
timestamp 1666464484
transform 1 0 36064 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1341_
timestamp 1666464484
transform 1 0 35052 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1342_
timestamp 1666464484
transform -1 0 36248 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1343_
timestamp 1666464484
transform 1 0 34960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1344_
timestamp 1666464484
transform 1 0 29716 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1345_
timestamp 1666464484
transform 1 0 34868 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1346_
timestamp 1666464484
transform 1 0 35512 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1347_
timestamp 1666464484
transform -1 0 40756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1348_
timestamp 1666464484
transform 1 0 39928 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _1349_
timestamp 1666464484
transform 1 0 40664 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1350_
timestamp 1666464484
transform 1 0 35788 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1351_
timestamp 1666464484
transform -1 0 37076 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1352_
timestamp 1666464484
transform -1 0 37812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1353_
timestamp 1666464484
transform 1 0 37628 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1354_
timestamp 1666464484
transform -1 0 34960 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1355_
timestamp 1666464484
transform -1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1356_
timestamp 1666464484
transform 1 0 40572 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_4  _1357_
timestamp 1666464484
transform 1 0 41308 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1666464484
transform 1 0 33672 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1359_
timestamp 1666464484
transform -1 0 34408 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1360_
timestamp 1666464484
transform -1 0 36892 0 1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_1  _1361_
timestamp 1666464484
transform 1 0 32292 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1362_
timestamp 1666464484
transform -1 0 32200 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _1363_
timestamp 1666464484
transform -1 0 34960 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__a31o_1  _1364_
timestamp 1666464484
transform 1 0 38180 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1365_
timestamp 1666464484
transform -1 0 39008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1366_
timestamp 1666464484
transform 1 0 38364 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1367_
timestamp 1666464484
transform 1 0 38824 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1368_
timestamp 1666464484
transform -1 0 39100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1369_
timestamp 1666464484
transform -1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1370_
timestamp 1666464484
transform -1 0 34224 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1371_
timestamp 1666464484
transform -1 0 36800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1372_
timestamp 1666464484
transform -1 0 36984 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1373_
timestamp 1666464484
transform 1 0 33856 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1374_
timestamp 1666464484
transform 1 0 33120 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1375_
timestamp 1666464484
transform 1 0 32752 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1376_
timestamp 1666464484
transform 1 0 32292 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1377_
timestamp 1666464484
transform -1 0 33212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_1  _1378_
timestamp 1666464484
transform 1 0 38824 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1379_
timestamp 1666464484
transform 1 0 39284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1380_
timestamp 1666464484
transform 1 0 39836 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1381_
timestamp 1666464484
transform -1 0 40572 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1382_
timestamp 1666464484
transform 1 0 38732 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1383_
timestamp 1666464484
transform -1 0 40664 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1384_
timestamp 1666464484
transform 1 0 40112 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1385_
timestamp 1666464484
transform 1 0 41216 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1386_
timestamp 1666464484
transform 1 0 41124 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1387_
timestamp 1666464484
transform -1 0 41492 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1388_
timestamp 1666464484
transform 1 0 41124 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1389_
timestamp 1666464484
transform 1 0 41768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1390_
timestamp 1666464484
transform -1 0 41768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1391_
timestamp 1666464484
transform 1 0 35328 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1392_
timestamp 1666464484
transform 1 0 40480 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1393_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 32384 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1394_
timestamp 1666464484
transform 1 0 41124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1395_
timestamp 1666464484
transform 1 0 41124 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _1396_
timestamp 1666464484
transform 1 0 34868 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1397_
timestamp 1666464484
transform -1 0 37904 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1398_
timestamp 1666464484
transform -1 0 35236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1399_
timestamp 1666464484
transform 1 0 33764 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _1400_
timestamp 1666464484
transform 1 0 35328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1401_
timestamp 1666464484
transform 1 0 34592 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1402_
timestamp 1666464484
transform 1 0 35052 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1403_
timestamp 1666464484
transform -1 0 35328 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1404_
timestamp 1666464484
transform 1 0 33396 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1405_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36064 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1406_
timestamp 1666464484
transform -1 0 38272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1666464484
transform 1 0 36432 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1408_
timestamp 1666464484
transform -1 0 37352 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1409_
timestamp 1666464484
transform -1 0 36984 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1410_
timestamp 1666464484
transform 1 0 37444 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1411_
timestamp 1666464484
transform 1 0 36708 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1412_
timestamp 1666464484
transform -1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1413_
timestamp 1666464484
transform 1 0 38180 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1414_
timestamp 1666464484
transform 1 0 37628 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1415_
timestamp 1666464484
transform 1 0 32108 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1416_
timestamp 1666464484
transform 1 0 36708 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1417_
timestamp 1666464484
transform 1 0 34960 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1418_
timestamp 1666464484
transform 1 0 36432 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1419_
timestamp 1666464484
transform -1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1420_
timestamp 1666464484
transform -1 0 37260 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1421_
timestamp 1666464484
transform 1 0 38640 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1422_
timestamp 1666464484
transform 1 0 40112 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1423_
timestamp 1666464484
transform 1 0 39928 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _1424_
timestamp 1666464484
transform -1 0 42228 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1425_
timestamp 1666464484
transform 1 0 42596 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1426_
timestamp 1666464484
transform -1 0 38088 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1427_
timestamp 1666464484
transform 1 0 38732 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1428_
timestamp 1666464484
transform -1 0 36800 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1429_
timestamp 1666464484
transform 1 0 36156 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1430_
timestamp 1666464484
transform -1 0 36616 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1431_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 36708 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1432_
timestamp 1666464484
transform 1 0 35696 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _1433_
timestamp 1666464484
transform 1 0 34868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1434_
timestamp 1666464484
transform 1 0 38548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1435_
timestamp 1666464484
transform 1 0 38364 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1436_
timestamp 1666464484
transform 1 0 37812 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1666464484
transform 1 0 37812 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1438_
timestamp 1666464484
transform 1 0 37444 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1439_
timestamp 1666464484
transform 1 0 38916 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1440_
timestamp 1666464484
transform 1 0 38456 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1441_
timestamp 1666464484
transform 1 0 38456 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1442_
timestamp 1666464484
transform -1 0 39560 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1443_
timestamp 1666464484
transform 1 0 39100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1444_
timestamp 1666464484
transform -1 0 40756 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1445_
timestamp 1666464484
transform 1 0 40020 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1446_
timestamp 1666464484
transform 1 0 41124 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1447_
timestamp 1666464484
transform 1 0 40480 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1448_
timestamp 1666464484
transform 1 0 40940 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1449_
timestamp 1666464484
transform 1 0 40112 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1450_
timestamp 1666464484
transform 1 0 39836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1451_
timestamp 1666464484
transform -1 0 37628 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1452_
timestamp 1666464484
transform 1 0 38180 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1453_
timestamp 1666464484
transform 1 0 33948 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1454_
timestamp 1666464484
transform 1 0 34868 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1455_
timestamp 1666464484
transform 1 0 37260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1666464484
transform -1 0 36248 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1457_
timestamp 1666464484
transform 1 0 35328 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1458_
timestamp 1666464484
transform 1 0 36432 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1459_
timestamp 1666464484
transform -1 0 36984 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1460_
timestamp 1666464484
transform -1 0 37812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_2  _1461_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36708 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1462_
timestamp 1666464484
transform 1 0 36064 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1463_
timestamp 1666464484
transform 1 0 35604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1464_
timestamp 1666464484
transform 1 0 37076 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1465_
timestamp 1666464484
transform -1 0 38640 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1466_
timestamp 1666464484
transform 1 0 39008 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1467_
timestamp 1666464484
transform -1 0 39192 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1468_
timestamp 1666464484
transform 1 0 40020 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1469_
timestamp 1666464484
transform 1 0 39928 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1470_
timestamp 1666464484
transform 1 0 40112 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1471_
timestamp 1666464484
transform 1 0 40020 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1472_
timestamp 1666464484
transform -1 0 41400 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1473_
timestamp 1666464484
transform 1 0 36616 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1474_
timestamp 1666464484
transform 1 0 37444 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1475_
timestamp 1666464484
transform -1 0 35604 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1476_
timestamp 1666464484
transform 1 0 34316 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1477_
timestamp 1666464484
transform -1 0 34960 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1478_
timestamp 1666464484
transform 1 0 34960 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1479_
timestamp 1666464484
transform 1 0 34132 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1480_
timestamp 1666464484
transform -1 0 36616 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1481_
timestamp 1666464484
transform 1 0 35880 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1482_
timestamp 1666464484
transform 1 0 37168 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1483_
timestamp 1666464484
transform 1 0 37444 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1484_
timestamp 1666464484
transform 1 0 37996 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1485_
timestamp 1666464484
transform 1 0 38456 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1486_
timestamp 1666464484
transform -1 0 40112 0 -1 26112
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1487_
timestamp 1666464484
transform -1 0 35972 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1488_
timestamp 1666464484
transform -1 0 35328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1489_
timestamp 1666464484
transform 1 0 35236 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1490_
timestamp 1666464484
transform 1 0 38364 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1491_
timestamp 1666464484
transform -1 0 39008 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1492_
timestamp 1666464484
transform -1 0 35420 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1493_
timestamp 1666464484
transform -1 0 39468 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1494_
timestamp 1666464484
transform -1 0 23920 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _1495_
timestamp 1666464484
transform 1 0 54832 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1496_
timestamp 1666464484
transform 1 0 53176 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1497_
timestamp 1666464484
transform 1 0 42596 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1498_
timestamp 1666464484
transform -1 0 53452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1499_
timestamp 1666464484
transform 1 0 41492 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  _1500_
timestamp 1666464484
transform 1 0 49312 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1501_
timestamp 1666464484
transform -1 0 52532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _1502_
timestamp 1666464484
transform 1 0 41400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1503_
timestamp 1666464484
transform -1 0 51704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1504_
timestamp 1666464484
transform -1 0 48116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1505_
timestamp 1666464484
transform -1 0 43700 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_2  _1506_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 54832 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 1666464484
transform -1 0 48024 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 1666464484
transform 1 0 44344 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1509_
timestamp 1666464484
transform 1 0 48116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1510_
timestamp 1666464484
transform -1 0 51428 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1511_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 50508 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1512_
timestamp 1666464484
transform 1 0 46828 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1513_
timestamp 1666464484
transform -1 0 48116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_2  _1514_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 50968 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1515_
timestamp 1666464484
transform -1 0 52440 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1516_
timestamp 1666464484
transform 1 0 43884 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1517_
timestamp 1666464484
transform -1 0 55936 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1518_
timestamp 1666464484
transform 1 0 50232 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1519_
timestamp 1666464484
transform -1 0 49864 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _1520_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 47012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _1521_
timestamp 1666464484
transform -1 0 56396 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_4  _1522_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 45356 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1523_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 44068 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1524_
timestamp 1666464484
transform -1 0 53728 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1525_
timestamp 1666464484
transform -1 0 49680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1526_
timestamp 1666464484
transform 1 0 43700 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1527_
timestamp 1666464484
transform 1 0 45908 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1528_
timestamp 1666464484
transform -1 0 47012 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _1529_
timestamp 1666464484
transform -1 0 55016 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_2  _1530_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 48024 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1531_
timestamp 1666464484
transform 1 0 48760 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1532_
timestamp 1666464484
transform 1 0 46092 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1533_
timestamp 1666464484
transform -1 0 43884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1534_
timestamp 1666464484
transform -1 0 44804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1535_
timestamp 1666464484
transform 1 0 42964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1536_
timestamp 1666464484
transform -1 0 45724 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1537_
timestamp 1666464484
transform 1 0 43608 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_4  _1538_
timestamp 1666464484
transform 1 0 42596 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__and2b_2  _1539_
timestamp 1666464484
transform -1 0 51060 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1540_
timestamp 1666464484
transform 1 0 50784 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1541_
timestamp 1666464484
transform 1 0 44620 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1542_
timestamp 1666464484
transform 1 0 44620 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_2  _1543_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 45540 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1544_
timestamp 1666464484
transform -1 0 45356 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _1545_
timestamp 1666464484
transform -1 0 48944 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _1546_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 48484 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__and3_1  _1547_
timestamp 1666464484
transform 1 0 48208 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1548_
timestamp 1666464484
transform 1 0 48944 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_2  _1549_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 54096 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1550_
timestamp 1666464484
transform -1 0 49404 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1551_
timestamp 1666464484
transform 1 0 48024 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1552_
timestamp 1666464484
transform -1 0 47748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1553_
timestamp 1666464484
transform 1 0 50324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1554_
timestamp 1666464484
transform 1 0 47288 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _1555_
timestamp 1666464484
transform -1 0 53176 0 1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_4  _1556_
timestamp 1666464484
transform 1 0 52348 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_2  _1557_
timestamp 1666464484
transform 1 0 54188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1558_
timestamp 1666464484
transform 1 0 46736 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1559_
timestamp 1666464484
transform 1 0 52624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1560_
timestamp 1666464484
transform 1 0 46460 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1561_
timestamp 1666464484
transform 1 0 44068 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1562_
timestamp 1666464484
transform 1 0 46828 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1563_
timestamp 1666464484
transform 1 0 47380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1564_
timestamp 1666464484
transform -1 0 43792 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1565_
timestamp 1666464484
transform -1 0 43424 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1566_
timestamp 1666464484
transform 1 0 43792 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1567_
timestamp 1666464484
transform -1 0 44528 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _1568_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43884 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _1569_
timestamp 1666464484
transform -1 0 45632 0 -1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1570_
timestamp 1666464484
transform 1 0 45816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1571_
timestamp 1666464484
transform 1 0 46828 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1572_
timestamp 1666464484
transform 1 0 48852 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _1573_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 55200 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _1574_
timestamp 1666464484
transform 1 0 49404 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1575_
timestamp 1666464484
transform 1 0 47840 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1576_
timestamp 1666464484
transform -1 0 46368 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1577_
timestamp 1666464484
transform 1 0 51520 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1578_
timestamp 1666464484
transform -1 0 52164 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1579_
timestamp 1666464484
transform -1 0 47104 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_2  _1580_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 45540 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1581_
timestamp 1666464484
transform 1 0 45264 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1582_
timestamp 1666464484
transform -1 0 55844 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1583_
timestamp 1666464484
transform -1 0 45540 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1584_
timestamp 1666464484
transform -1 0 51336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1585_
timestamp 1666464484
transform 1 0 48668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1586_
timestamp 1666464484
transform 1 0 49864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1587_
timestamp 1666464484
transform 1 0 44252 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1588_
timestamp 1666464484
transform 1 0 49404 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1589_
timestamp 1666464484
transform -1 0 54004 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1590_
timestamp 1666464484
transform -1 0 51980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1591_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 50692 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _1592_
timestamp 1666464484
transform -1 0 53544 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1593_
timestamp 1666464484
transform 1 0 48760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1594_
timestamp 1666464484
transform 1 0 49036 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1595_
timestamp 1666464484
transform -1 0 48300 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1596_
timestamp 1666464484
transform 1 0 47656 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1597_
timestamp 1666464484
transform -1 0 46552 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1598_
timestamp 1666464484
transform -1 0 46276 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1599_
timestamp 1666464484
transform -1 0 47104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1600_
timestamp 1666464484
transform 1 0 52900 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1601_
timestamp 1666464484
transform -1 0 48668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1602_
timestamp 1666464484
transform -1 0 43148 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _1603_
timestamp 1666464484
transform -1 0 43792 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1604_
timestamp 1666464484
transform -1 0 45632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1605_
timestamp 1666464484
transform -1 0 44068 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1606_
timestamp 1666464484
transform 1 0 46368 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1607_
timestamp 1666464484
transform 1 0 45172 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1608_
timestamp 1666464484
transform -1 0 47840 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1609_
timestamp 1666464484
transform -1 0 48116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1610_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 46368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1611_
timestamp 1666464484
transform -1 0 48300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1612_
timestamp 1666464484
transform -1 0 47012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1613_
timestamp 1666464484
transform -1 0 49864 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1614_
timestamp 1666464484
transform 1 0 51244 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1615_
timestamp 1666464484
transform -1 0 50876 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1616_
timestamp 1666464484
transform -1 0 51888 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1617_
timestamp 1666464484
transform 1 0 49128 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1618_
timestamp 1666464484
transform 1 0 48944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1619_
timestamp 1666464484
transform -1 0 49680 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1620_
timestamp 1666464484
transform -1 0 44528 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1621_
timestamp 1666464484
transform 1 0 44252 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _1622_
timestamp 1666464484
transform 1 0 45540 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1623_
timestamp 1666464484
transform -1 0 48024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1624_
timestamp 1666464484
transform -1 0 47380 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _1625_
timestamp 1666464484
transform 1 0 45724 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1626_
timestamp 1666464484
transform 1 0 46000 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1627_
timestamp 1666464484
transform 1 0 55476 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1628_
timestamp 1666464484
transform 1 0 45356 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1629_
timestamp 1666464484
transform 1 0 41768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1630_
timestamp 1666464484
transform 1 0 45172 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1631_
timestamp 1666464484
transform 1 0 44252 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _1632_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 42044 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1633_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 42964 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1634_
timestamp 1666464484
transform 1 0 45172 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1635_
timestamp 1666464484
transform 1 0 43792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_1  _1636_
timestamp 1666464484
transform -1 0 46184 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1637_
timestamp 1666464484
transform -1 0 45356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1638_
timestamp 1666464484
transform 1 0 43976 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1639_
timestamp 1666464484
transform -1 0 43700 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1640_
timestamp 1666464484
transform -1 0 44528 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1641_
timestamp 1666464484
transform -1 0 44252 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1642_
timestamp 1666464484
transform 1 0 43056 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _1643_
timestamp 1666464484
transform -1 0 44620 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1644_
timestamp 1666464484
transform -1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1645_
timestamp 1666464484
transform 1 0 44068 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1646_
timestamp 1666464484
transform 1 0 46736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1647_
timestamp 1666464484
transform 1 0 45816 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _1648_
timestamp 1666464484
transform -1 0 43884 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1649_
timestamp 1666464484
transform -1 0 46736 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1650_
timestamp 1666464484
transform -1 0 45724 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1651_
timestamp 1666464484
transform 1 0 46460 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1652_
timestamp 1666464484
transform -1 0 46276 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _1653_
timestamp 1666464484
transform -1 0 45816 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1654_
timestamp 1666464484
transform 1 0 45356 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1655_
timestamp 1666464484
transform -1 0 45632 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1656_
timestamp 1666464484
transform -1 0 43976 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1657_
timestamp 1666464484
transform 1 0 43516 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _1658_
timestamp 1666464484
transform 1 0 45172 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1659_
timestamp 1666464484
transform -1 0 46828 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1660_
timestamp 1666464484
transform 1 0 45908 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1661_
timestamp 1666464484
transform 1 0 47196 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1662_
timestamp 1666464484
transform -1 0 47104 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1663_
timestamp 1666464484
transform 1 0 44160 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_4  _1664_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 44160 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__and2b_1  _1665_
timestamp 1666464484
transform 1 0 44804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1666_
timestamp 1666464484
transform -1 0 47748 0 1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__and3_1  _1667_
timestamp 1666464484
transform 1 0 45724 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1668_
timestamp 1666464484
transform 1 0 46368 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1669_
timestamp 1666464484
transform 1 0 46736 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1670_
timestamp 1666464484
transform -1 0 47748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1671_
timestamp 1666464484
transform 1 0 47748 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1672_
timestamp 1666464484
transform 1 0 46000 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1673_
timestamp 1666464484
transform -1 0 41676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1674_
timestamp 1666464484
transform 1 0 42044 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1675_
timestamp 1666464484
transform -1 0 46000 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1676_
timestamp 1666464484
transform 1 0 46552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1677_
timestamp 1666464484
transform 1 0 46920 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1678_
timestamp 1666464484
transform 1 0 47380 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1679_
timestamp 1666464484
transform 1 0 45632 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1680_
timestamp 1666464484
transform 1 0 46460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1681_
timestamp 1666464484
transform 1 0 42688 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1682_
timestamp 1666464484
transform -1 0 43056 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1683_
timestamp 1666464484
transform -1 0 47932 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1684_
timestamp 1666464484
transform 1 0 47748 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1685_
timestamp 1666464484
transform 1 0 48484 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _1686_
timestamp 1666464484
transform -1 0 48576 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1687_
timestamp 1666464484
transform -1 0 48208 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1688_
timestamp 1666464484
transform 1 0 46920 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _1689_
timestamp 1666464484
transform -1 0 48208 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1690_
timestamp 1666464484
transform -1 0 48392 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1691_
timestamp 1666464484
transform -1 0 47288 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1692_
timestamp 1666464484
transform -1 0 54648 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _1693_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 53544 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1694_
timestamp 1666464484
transform 1 0 51888 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1695_
timestamp 1666464484
transform 1 0 54648 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1696_
timestamp 1666464484
transform -1 0 51152 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1697_
timestamp 1666464484
transform -1 0 50876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1698_
timestamp 1666464484
transform 1 0 51704 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1699_
timestamp 1666464484
transform 1 0 50600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1700_
timestamp 1666464484
transform -1 0 50876 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1701_
timestamp 1666464484
transform 1 0 44252 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1702_
timestamp 1666464484
transform -1 0 48208 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1703_
timestamp 1666464484
transform 1 0 47012 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1704_
timestamp 1666464484
transform 1 0 47656 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1705_
timestamp 1666464484
transform 1 0 46736 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1706_
timestamp 1666464484
transform 1 0 47840 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1707_
timestamp 1666464484
transform 1 0 47932 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1708_
timestamp 1666464484
transform -1 0 49312 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _1709_
timestamp 1666464484
transform -1 0 46736 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1710_
timestamp 1666464484
transform 1 0 48116 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1711_
timestamp 1666464484
transform 1 0 44436 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1712_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 45448 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1713_
timestamp 1666464484
transform -1 0 42596 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1714_
timestamp 1666464484
transform 1 0 41400 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1715_
timestamp 1666464484
transform 1 0 45632 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1716_
timestamp 1666464484
transform -1 0 42872 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1717_
timestamp 1666464484
transform 1 0 45172 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1718_
timestamp 1666464484
transform -1 0 46276 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1719_
timestamp 1666464484
transform 1 0 47564 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1720_
timestamp 1666464484
transform 1 0 48024 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1721_
timestamp 1666464484
transform 1 0 53084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1722_
timestamp 1666464484
transform 1 0 53728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1723_
timestamp 1666464484
transform 1 0 55476 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1724_
timestamp 1666464484
transform 1 0 56304 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1725_
timestamp 1666464484
transform -1 0 54464 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1726_
timestamp 1666464484
transform 1 0 51244 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1727_
timestamp 1666464484
transform -1 0 51060 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1728_
timestamp 1666464484
transform -1 0 50784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1729_
timestamp 1666464484
transform -1 0 51796 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _1730_
timestamp 1666464484
transform -1 0 49220 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1731_
timestamp 1666464484
transform -1 0 49404 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1732_
timestamp 1666464484
transform -1 0 48944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1733_
timestamp 1666464484
transform -1 0 48392 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1734_
timestamp 1666464484
transform 1 0 48300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1735_
timestamp 1666464484
transform -1 0 48944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1736_
timestamp 1666464484
transform 1 0 48300 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1737_
timestamp 1666464484
transform 1 0 49404 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _1738_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 49404 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1739_
timestamp 1666464484
transform -1 0 49588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1740_
timestamp 1666464484
transform 1 0 48852 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1741_
timestamp 1666464484
transform -1 0 49036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1742_
timestamp 1666464484
transform 1 0 48576 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1743_
timestamp 1666464484
transform 1 0 49680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1744_
timestamp 1666464484
transform 1 0 48944 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1745_
timestamp 1666464484
transform 1 0 43700 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1746_
timestamp 1666464484
transform 1 0 48300 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1747_
timestamp 1666464484
transform 1 0 43240 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1748_
timestamp 1666464484
transform 1 0 43516 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1749_
timestamp 1666464484
transform 1 0 48024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1750_
timestamp 1666464484
transform -1 0 49312 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1751_
timestamp 1666464484
transform 1 0 49312 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1752_
timestamp 1666464484
transform 1 0 48300 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1753_
timestamp 1666464484
transform 1 0 49128 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _1754_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 48760 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o21bai_2  _1755_
timestamp 1666464484
transform -1 0 48576 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_4  _1756_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 49312 0 -1 28288
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_1  _1757_
timestamp 1666464484
transform 1 0 49220 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_4  _1758_
timestamp 1666464484
transform -1 0 51060 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1759_
timestamp 1666464484
transform -1 0 49864 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1760_
timestamp 1666464484
transform 1 0 49220 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1761_
timestamp 1666464484
transform -1 0 50784 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1762_
timestamp 1666464484
transform 1 0 41860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1763_
timestamp 1666464484
transform 1 0 49680 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1764_
timestamp 1666464484
transform 1 0 46092 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1765_
timestamp 1666464484
transform -1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1766_
timestamp 1666464484
transform 1 0 45724 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1767_
timestamp 1666464484
transform -1 0 46460 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1768_
timestamp 1666464484
transform -1 0 50416 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1769_
timestamp 1666464484
transform 1 0 49496 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1770_
timestamp 1666464484
transform 1 0 46736 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a311o_1  _1771_
timestamp 1666464484
transform -1 0 47104 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1772_
timestamp 1666464484
transform -1 0 47196 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1773_
timestamp 1666464484
transform 1 0 46552 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1774_
timestamp 1666464484
transform 1 0 47748 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1775_
timestamp 1666464484
transform 1 0 48760 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1776_
timestamp 1666464484
transform 1 0 48852 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1777_
timestamp 1666464484
transform -1 0 49864 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1778_
timestamp 1666464484
transform -1 0 49956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1779_
timestamp 1666464484
transform 1 0 50140 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1780_
timestamp 1666464484
transform 1 0 48760 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1781_
timestamp 1666464484
transform 1 0 50416 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1782_
timestamp 1666464484
transform -1 0 52440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1783_
timestamp 1666464484
transform 1 0 52808 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1784_
timestamp 1666464484
transform -1 0 52440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1785_
timestamp 1666464484
transform 1 0 54740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1786_
timestamp 1666464484
transform -1 0 50692 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1787_
timestamp 1666464484
transform 1 0 55476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1788_
timestamp 1666464484
transform 1 0 52992 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1789_
timestamp 1666464484
transform 1 0 51888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1790_
timestamp 1666464484
transform -1 0 51060 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1791_
timestamp 1666464484
transform 1 0 50324 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1792_
timestamp 1666464484
transform -1 0 50968 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1793_
timestamp 1666464484
transform 1 0 50784 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1794_
timestamp 1666464484
transform 1 0 51428 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1795_
timestamp 1666464484
transform 1 0 50784 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1796_
timestamp 1666464484
transform 1 0 51428 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1797_
timestamp 1666464484
transform -1 0 51152 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1798_
timestamp 1666464484
transform -1 0 54372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1799_
timestamp 1666464484
transform 1 0 55476 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1800_
timestamp 1666464484
transform 1 0 55568 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1801_
timestamp 1666464484
transform 1 0 55476 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _1802_
timestamp 1666464484
transform -1 0 53452 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1803_
timestamp 1666464484
transform 1 0 51796 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1804_
timestamp 1666464484
transform -1 0 48392 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1805_
timestamp 1666464484
transform 1 0 51520 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1806_
timestamp 1666464484
transform 1 0 44528 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1807_
timestamp 1666464484
transform -1 0 43976 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1808_
timestamp 1666464484
transform 1 0 42688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1809_
timestamp 1666464484
transform 1 0 43424 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1810_
timestamp 1666464484
transform -1 0 43976 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1811_
timestamp 1666464484
transform 1 0 45632 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1812_
timestamp 1666464484
transform 1 0 50416 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1813_
timestamp 1666464484
transform -1 0 52440 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1814_
timestamp 1666464484
transform 1 0 51888 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1815_
timestamp 1666464484
transform 1 0 52900 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1816_
timestamp 1666464484
transform 1 0 51244 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1817_
timestamp 1666464484
transform -1 0 56120 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _1818_
timestamp 1666464484
transform 1 0 50784 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1819_
timestamp 1666464484
transform -1 0 51336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1820_
timestamp 1666464484
transform -1 0 52624 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1821_
timestamp 1666464484
transform 1 0 51612 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1822_
timestamp 1666464484
transform -1 0 53268 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_2  _1823_
timestamp 1666464484
transform 1 0 50324 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _1824_
timestamp 1666464484
transform 1 0 51888 0 1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__a311oi_4  _1825_
timestamp 1666464484
transform 1 0 51152 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__a31o_1  _1826_
timestamp 1666464484
transform -1 0 51612 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1827_
timestamp 1666464484
transform 1 0 52164 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1828_
timestamp 1666464484
transform 1 0 52900 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1829_
timestamp 1666464484
transform 1 0 58052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1830_
timestamp 1666464484
transform 1 0 54372 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1831_
timestamp 1666464484
transform 1 0 53636 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1832_
timestamp 1666464484
transform 1 0 54004 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1833_
timestamp 1666464484
transform 1 0 53820 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1834_
timestamp 1666464484
transform 1 0 54280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1835_
timestamp 1666464484
transform -1 0 52900 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1836_
timestamp 1666464484
transform 1 0 49404 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1837_
timestamp 1666464484
transform -1 0 50876 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1838_
timestamp 1666464484
transform 1 0 52072 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1839_
timestamp 1666464484
transform -1 0 53268 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1840_
timestamp 1666464484
transform 1 0 52900 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1841_
timestamp 1666464484
transform 1 0 51704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1842_
timestamp 1666464484
transform 1 0 50140 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1843_
timestamp 1666464484
transform -1 0 50692 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1844_
timestamp 1666464484
transform 1 0 50324 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1845_
timestamp 1666464484
transform 1 0 53268 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _1846_
timestamp 1666464484
transform 1 0 53360 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1847_
timestamp 1666464484
transform 1 0 53360 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1848_
timestamp 1666464484
transform 1 0 53636 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1849_
timestamp 1666464484
transform -1 0 53268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1850_
timestamp 1666464484
transform 1 0 54004 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1851_
timestamp 1666464484
transform 1 0 53544 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1852_
timestamp 1666464484
transform 1 0 53636 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1853_
timestamp 1666464484
transform -1 0 52440 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1854_
timestamp 1666464484
transform -1 0 53452 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1855_
timestamp 1666464484
transform -1 0 55200 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1856_
timestamp 1666464484
transform 1 0 53912 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1857_
timestamp 1666464484
transform 1 0 53912 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1858_
timestamp 1666464484
transform 1 0 52164 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1859_
timestamp 1666464484
transform 1 0 54556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1860_
timestamp 1666464484
transform 1 0 53544 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1861_
timestamp 1666464484
transform -1 0 55016 0 1 26112
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1862_
timestamp 1666464484
transform -1 0 52440 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1863_
timestamp 1666464484
transform -1 0 53452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1864_
timestamp 1666464484
transform -1 0 52992 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1865_
timestamp 1666464484
transform -1 0 51704 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1866_
timestamp 1666464484
transform -1 0 51888 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1867_
timestamp 1666464484
transform -1 0 54004 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1868_
timestamp 1666464484
transform 1 0 51336 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1869_
timestamp 1666464484
transform 1 0 50048 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_2  _1870_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 50876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1871_
timestamp 1666464484
transform 1 0 43516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1872_
timestamp 1666464484
transform -1 0 52900 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1873_
timestamp 1666464484
transform 1 0 52992 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1874_
timestamp 1666464484
transform 1 0 53820 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _1875_
timestamp 1666464484
transform 1 0 54096 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1876_
timestamp 1666464484
transform 1 0 54096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _1877_
timestamp 1666464484
transform 1 0 54648 0 -1 25024
box -38 -48 2062 592
use sky130_fd_sc_hd__a221oi_4  _1878_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 50508 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _1879_
timestamp 1666464484
transform 1 0 55016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1880_
timestamp 1666464484
transform -1 0 56120 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1881_
timestamp 1666464484
transform -1 0 56212 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _1882_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 55016 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _1883_
timestamp 1666464484
transform -1 0 57500 0 1 26112
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _1884_
timestamp 1666464484
transform -1 0 53268 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1885_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 53820 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1886_
timestamp 1666464484
transform -1 0 57224 0 -1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _1887_
timestamp 1666464484
transform 1 0 54280 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1888_
timestamp 1666464484
transform -1 0 54188 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1889_
timestamp 1666464484
transform -1 0 55016 0 -1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _1890_
timestamp 1666464484
transform 1 0 55476 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1891_
timestamp 1666464484
transform 1 0 55200 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1892_
timestamp 1666464484
transform -1 0 53636 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1893_
timestamp 1666464484
transform -1 0 53820 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1894_
timestamp 1666464484
transform 1 0 53820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1895_
timestamp 1666464484
transform -1 0 54004 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1896_
timestamp 1666464484
transform 1 0 51612 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1897_
timestamp 1666464484
transform -1 0 51704 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1898_
timestamp 1666464484
transform 1 0 54464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1899_
timestamp 1666464484
transform -1 0 54924 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1900_
timestamp 1666464484
transform 1 0 53912 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1901_
timestamp 1666464484
transform -1 0 54648 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1902_
timestamp 1666464484
transform 1 0 55016 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1903_
timestamp 1666464484
transform 1 0 55476 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1904_
timestamp 1666464484
transform 1 0 54924 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1905_
timestamp 1666464484
transform -1 0 56212 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1906_
timestamp 1666464484
transform -1 0 56856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1907_
timestamp 1666464484
transform 1 0 55476 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1908_
timestamp 1666464484
transform 1 0 55476 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1909_
timestamp 1666464484
transform 1 0 55844 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1910_
timestamp 1666464484
transform 1 0 56028 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1911_
timestamp 1666464484
transform -1 0 58328 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1912_
timestamp 1666464484
transform 1 0 55844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1666464484
transform 1 0 55476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o311ai_4  _1914_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 52900 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _1915_
timestamp 1666464484
transform 1 0 56764 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _1916_
timestamp 1666464484
transform -1 0 58420 0 1 27200
box -38 -48 2062 592
use sky130_fd_sc_hd__or2b_1  _1917_
timestamp 1666464484
transform 1 0 55568 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1918_
timestamp 1666464484
transform 1 0 51980 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1919_
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1920_
timestamp 1666464484
transform 1 0 50968 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1921_
timestamp 1666464484
transform 1 0 52900 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1922_
timestamp 1666464484
transform -1 0 53544 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1923_
timestamp 1666464484
transform 1 0 52900 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1924_
timestamp 1666464484
transform -1 0 53452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1925_
timestamp 1666464484
transform -1 0 53728 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1926_
timestamp 1666464484
transform 1 0 55476 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1927_
timestamp 1666464484
transform -1 0 56488 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1928_
timestamp 1666464484
transform -1 0 56856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1929_
timestamp 1666464484
transform 1 0 56488 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1930_
timestamp 1666464484
transform 1 0 56856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1931_
timestamp 1666464484
transform -1 0 56856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1932_
timestamp 1666464484
transform 1 0 56580 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1933_
timestamp 1666464484
transform 1 0 57224 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1934_
timestamp 1666464484
transform 1 0 58052 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1935_
timestamp 1666464484
transform -1 0 57592 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1936_
timestamp 1666464484
transform -1 0 58420 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _1937_
timestamp 1666464484
transform 1 0 55568 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1938_
timestamp 1666464484
transform -1 0 51060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1939_
timestamp 1666464484
transform -1 0 51152 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_2  _1940_
timestamp 1666464484
transform 1 0 50416 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1941_
timestamp 1666464484
transform 1 0 56580 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1942_
timestamp 1666464484
transform 1 0 57316 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1943_
timestamp 1666464484
transform -1 0 58420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1944_
timestamp 1666464484
transform 1 0 57500 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1945_
timestamp 1666464484
transform 1 0 58052 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1946_
timestamp 1666464484
transform 1 0 56856 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1947_
timestamp 1666464484
transform 1 0 57040 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1948_
timestamp 1666464484
transform 1 0 57684 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1949_
timestamp 1666464484
transform 1 0 52440 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1950_
timestamp 1666464484
transform 1 0 56212 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1951_
timestamp 1666464484
transform -1 0 55844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1952_
timestamp 1666464484
transform -1 0 56580 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1953_
timestamp 1666464484
transform -1 0 58328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1954_
timestamp 1666464484
transform 1 0 57592 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1955_
timestamp 1666464484
transform -1 0 57316 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1956_
timestamp 1666464484
transform -1 0 57224 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1957_
timestamp 1666464484
transform -1 0 46276 0 -1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  _1958_
timestamp 1666464484
transform 1 0 50324 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1959_
timestamp 1666464484
transform 1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1960_
timestamp 1666464484
transform 1 0 41032 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1961_
timestamp 1666464484
transform 1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1962_
timestamp 1666464484
transform -1 0 55200 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1963_
timestamp 1666464484
transform 1 0 41308 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1964_
timestamp 1666464484
transform -1 0 38732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1965_
timestamp 1666464484
transform 1 0 42412 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1966_
timestamp 1666464484
transform -1 0 39284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1967_
timestamp 1666464484
transform 1 0 40204 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1968_
timestamp 1666464484
transform 1 0 41032 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1969_
timestamp 1666464484
transform 1 0 42596 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1970_
timestamp 1666464484
transform 1 0 40940 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1971_
timestamp 1666464484
transform -1 0 42872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1972_
timestamp 1666464484
transform -1 0 43516 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1973_
timestamp 1666464484
transform -1 0 44344 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1974_
timestamp 1666464484
transform 1 0 43976 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _1975_
timestamp 1666464484
transform -1 0 45724 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1976_
timestamp 1666464484
transform 1 0 45448 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1977_
timestamp 1666464484
transform 1 0 46092 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1978_
timestamp 1666464484
transform -1 0 40664 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1979_
timestamp 1666464484
transform -1 0 37628 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1980_
timestamp 1666464484
transform 1 0 39284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1981_
timestamp 1666464484
transform -1 0 38180 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1982_
timestamp 1666464484
transform -1 0 39192 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1983_
timestamp 1666464484
transform -1 0 39376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1984_
timestamp 1666464484
transform -1 0 38732 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1985_
timestamp 1666464484
transform -1 0 41216 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1986_
timestamp 1666464484
transform 1 0 41032 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1987_
timestamp 1666464484
transform -1 0 40848 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1988_
timestamp 1666464484
transform -1 0 40664 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1989_
timestamp 1666464484
transform -1 0 23368 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1990_
timestamp 1666464484
transform -1 0 22264 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1991_
timestamp 1666464484
transform -1 0 53360 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1992_
timestamp 1666464484
transform 1 0 47748 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1993_
timestamp 1666464484
transform 1 0 47012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1994_
timestamp 1666464484
transform 1 0 45172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1995_
timestamp 1666464484
transform -1 0 42872 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1996_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 45724 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1997_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1998_
timestamp 1666464484
transform 1 0 39744 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1999_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 45080 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2000_
timestamp 1666464484
transform -1 0 40664 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2001_
timestamp 1666464484
transform 1 0 37444 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2002_
timestamp 1666464484
transform -1 0 37904 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2003_
timestamp 1666464484
transform 1 0 42596 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2004_
timestamp 1666464484
transform -1 0 45356 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2005_
timestamp 1666464484
transform 1 0 38732 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2006_
timestamp 1666464484
transform -1 0 36984 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2007_
timestamp 1666464484
transform -1 0 35696 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2008_
timestamp 1666464484
transform 1 0 40940 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2009_
timestamp 1666464484
transform -1 0 44712 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2010_
timestamp 1666464484
transform -1 0 37720 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2011_
timestamp 1666464484
transform 1 0 21988 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2012_
timestamp 1666464484
transform 1 0 21988 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2013_
timestamp 1666464484
transform 1 0 44528 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dlxtn_1  _2014_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 42780 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _2015_
timestamp 1666464484
transform 1 0 42872 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2016_
timestamp 1666464484
transform 1 0 45816 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2017_
timestamp 1666464484
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _2018_
timestamp 1666464484
transform 1 0 23000 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _2019_
timestamp 1666464484
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2020_
timestamp 1666464484
transform 1 0 41676 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2021_
timestamp 1666464484
transform 1 0 42596 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 42044 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_CLK
timestamp 1666464484
transform -1 0 39284 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_CLK
timestamp 1666464484
transform 1 0 42596 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1666464484
transform 1 0 53268 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1666464484
transform 1 0 40020 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1666464484
transform -1 0 35236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1666464484
transform 1 0 43332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1666464484
transform -1 0 35604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1666464484
transform 1 0 43424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1666464484
transform 1 0 34868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1666464484
transform 1 0 22356 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1666464484
transform 1 0 1564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1666464484
transform 1 0 32292 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 6072 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1666464484
transform -1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1666464484
transform -1 0 56488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1666464484
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1666464484
transform 1 0 58052 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1666464484
transform -1 0 4324 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1666464484
transform -1 0 1932 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1666464484
transform -1 0 49404 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1666464484
transform -1 0 36340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1666464484
transform 1 0 58052 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1666464484
transform 1 0 58052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1666464484
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1666464484
transform -1 0 1932 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1666464484
transform -1 0 1932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1666464484
transform 1 0 38088 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1666464484
transform 1 0 55476 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1666464484
transform -1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1666464484
transform 1 0 58052 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1666464484
transform -1 0 15916 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666464484
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1666464484
transform -1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1666464484
transform 1 0 58052 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1666464484
transform -1 0 10120 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1666464484
transform -1 0 1932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1666464484
transform -1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666464484
transform -1 0 43608 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1666464484
transform 1 0 58052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1666464484
transform -1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1666464484
transform -1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1666464484
transform 1 0 58052 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1666464484
transform -1 0 28152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1666464484
transform 1 0 58052 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1666464484
transform 1 0 58052 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1666464484
transform -1 0 22356 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1666464484
transform -1 0 27508 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1666464484
transform 1 0 40020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1666464484
transform -1 0 1932 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1666464484
transform -1 0 1932 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1666464484
transform 1 0 58052 0 -1 25024
box -38 -48 406 592
<< labels >>
flabel metal3 s 200 17688 800 17808 0 FreeSans 480 0 0 0 BitIn
port 0 nsew signal input
flabel metal2 s 44454 200 44510 800 0 FreeSans 224 90 0 0 CLK
port 1 nsew signal input
flabel metal2 s 32218 59200 32274 59800 0 FreeSans 224 90 0 0 EN
port 2 nsew signal input
flabel metal3 s 200 46928 800 47048 0 FreeSans 480 0 0 0 I[0]
port 3 nsew signal tristate
flabel metal2 s 56046 200 56102 800 0 FreeSans 224 90 0 0 I[10]
port 4 nsew signal tristate
flabel metal3 s 59200 688 59800 808 0 FreeSans 480 0 0 0 I[11]
port 5 nsew signal tristate
flabel metal3 s 59200 36728 59800 36848 0 FreeSans 480 0 0 0 I[12]
port 6 nsew signal tristate
flabel metal2 s 3882 59200 3938 59800 0 FreeSans 224 90 0 0 I[1]
port 7 nsew signal tristate
flabel metal3 s 200 53048 800 53168 0 FreeSans 480 0 0 0 I[2]
port 8 nsew signal tristate
flabel metal2 s 48962 59200 49018 59800 0 FreeSans 224 90 0 0 I[3]
port 9 nsew signal tristate
flabel metal2 s 33506 200 33562 800 0 FreeSans 224 90 0 0 I[4]
port 10 nsew signal tristate
flabel metal3 s 59200 42168 59800 42288 0 FreeSans 480 0 0 0 I[5]
port 11 nsew signal tristate
flabel metal3 s 59200 6808 59800 6928 0 FreeSans 480 0 0 0 I[6]
port 12 nsew signal tristate
flabel metal2 s 10966 200 11022 800 0 FreeSans 224 90 0 0 I[7]
port 13 nsew signal tristate
flabel metal3 s 200 40808 800 40928 0 FreeSans 480 0 0 0 I[8]
port 14 nsew signal tristate
flabel metal3 s 200 29248 800 29368 0 FreeSans 480 0 0 0 I[9]
port 15 nsew signal tristate
flabel metal2 s 38014 59200 38070 59800 0 FreeSans 224 90 0 0 Q[0]
port 16 nsew signal tristate
flabel metal2 s 54758 59200 54814 59800 0 FreeSans 224 90 0 0 Q[10]
port 17 nsew signal tristate
flabel metal3 s 200 35368 800 35488 0 FreeSans 480 0 0 0 Q[11]
port 18 nsew signal tristate
flabel metal3 s 59200 48288 59800 48408 0 FreeSans 480 0 0 0 Q[12]
port 19 nsew signal tristate
flabel metal2 s 15474 59200 15530 59800 0 FreeSans 224 90 0 0 Q[1]
port 20 nsew signal tristate
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 Q[2]
port 21 nsew signal tristate
flabel metal3 s 200 11568 800 11688 0 FreeSans 480 0 0 0 Q[3]
port 22 nsew signal tristate
flabel metal3 s 59200 30608 59800 30728 0 FreeSans 480 0 0 0 Q[4]
port 23 nsew signal tristate
flabel metal2 s 9678 59200 9734 59800 0 FreeSans 224 90 0 0 Q[5]
port 24 nsew signal tristate
flabel metal3 s 200 5448 800 5568 0 FreeSans 480 0 0 0 Q[6]
port 25 nsew signal tristate
flabel metal2 s 50250 200 50306 800 0 FreeSans 224 90 0 0 Q[7]
port 26 nsew signal tristate
flabel metal2 s 43166 59200 43222 59800 0 FreeSans 224 90 0 0 Q[8]
port 27 nsew signal tristate
flabel metal3 s 59200 12928 59800 13048 0 FreeSans 480 0 0 0 Q[9]
port 28 nsew signal tristate
flabel metal2 s 5170 200 5226 800 0 FreeSans 224 90 0 0 RST
port 29 nsew signal input
flabel metal2 s 16762 200 16818 800 0 FreeSans 224 90 0 0 addI[0]
port 30 nsew signal tristate
flabel metal2 s 21914 200 21970 800 0 FreeSans 224 90 0 0 addI[1]
port 31 nsew signal tristate
flabel metal3 s 59200 18368 59800 18488 0 FreeSans 480 0 0 0 addI[2]
port 32 nsew signal tristate
flabel metal2 s 27710 200 27766 800 0 FreeSans 224 90 0 0 addI[3]
port 33 nsew signal tristate
flabel metal3 s 59200 54408 59800 54528 0 FreeSans 480 0 0 0 addI[4]
port 34 nsew signal tristate
flabel metal3 s 59200 59848 59800 59968 0 FreeSans 480 0 0 0 addI[5]
port 35 nsew signal tristate
flabel metal2 s 21270 59200 21326 59800 0 FreeSans 224 90 0 0 addQ[0]
port 36 nsew signal tristate
flabel metal2 s 26422 59200 26478 59800 0 FreeSans 224 90 0 0 addQ[1]
port 37 nsew signal tristate
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 addQ[2]
port 38 nsew signal tristate
flabel metal3 s 200 23128 800 23248 0 FreeSans 480 0 0 0 addQ[3]
port 39 nsew signal tristate
flabel metal3 s 200 59168 800 59288 0 FreeSans 480 0 0 0 addQ[4]
port 40 nsew signal tristate
flabel metal3 s 59200 24488 59800 24608 0 FreeSans 480 0 0 0 addQ[5]
port 41 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 42 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 42 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 43 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 43 nsew ground bidirectional
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel via2 1610 17765 1610 17765 0 BitIn
rlabel metal1 41998 4624 41998 4624 0 CLK
rlabel metal1 32292 57426 32292 57426 0 EN
rlabel metal3 1188 46988 1188 46988 0 I[0]
rlabel metal2 56074 1520 56074 1520 0 I[10]
rlabel metal1 59110 2278 59110 2278 0 I[11]
rlabel metal2 58282 36941 58282 36941 0 I[12]
rlabel metal1 4002 57562 4002 57562 0 I[1]
rlabel metal3 1188 53108 1188 53108 0 I[2]
rlabel metal1 49082 57562 49082 57562 0 I[3]
rlabel metal2 33534 1554 33534 1554 0 I[4]
rlabel metal2 58282 42381 58282 42381 0 I[5]
rlabel metal1 58098 7174 58098 7174 0 I[6]
rlabel metal2 10994 1520 10994 1520 0 I[7]
rlabel metal3 1188 40868 1188 40868 0 I[8]
rlabel metal3 1188 29308 1188 29308 0 I[9]
rlabel metal1 38180 57562 38180 57562 0 Q[0]
rlabel metal2 54786 58388 54786 58388 0 Q[10]
rlabel metal3 1188 35428 1188 35428 0 Q[11]
rlabel metal2 58282 48433 58282 48433 0 Q[12]
rlabel metal1 15594 57562 15594 57562 0 Q[1]
rlabel metal2 46 1520 46 1520 0 Q[2]
rlabel metal3 1188 11628 1188 11628 0 Q[3]
rlabel metal2 58282 30617 58282 30617 0 Q[4]
rlabel metal1 9798 57562 9798 57562 0 Q[5]
rlabel metal3 1188 5508 1188 5508 0 Q[6]
rlabel metal2 50278 1027 50278 1027 0 Q[7]
rlabel metal1 43286 57562 43286 57562 0 Q[8]
rlabel metal2 58282 13073 58282 13073 0 Q[9]
rlabel metal1 5796 2414 5796 2414 0 RST
rlabel metal2 41814 4216 41814 4216 0 Reg_Delay_Q.In
rlabel metal1 45770 2550 45770 2550 0 Reg_Delay_Q.Out
rlabel metal1 42964 19482 42964 19482 0 _0000_
rlabel metal2 42826 20060 42826 20060 0 _0001_
rlabel metal2 23322 14858 23322 14858 0 _0002_
rlabel metal1 23046 14484 23046 14484 0 _0003_
rlabel metal2 55246 15079 55246 15079 0 _0004_
rlabel metal1 22034 18292 22034 18292 0 _0005_
rlabel metal2 46874 5848 46874 5848 0 _0006_
rlabel metal1 38962 3638 38962 3638 0 _0007_
rlabel metal1 39376 3706 39376 3706 0 _0008_
rlabel metal2 45402 4964 45402 4964 0 _0009_
rlabel metal1 40710 5270 40710 5270 0 _0010_
rlabel metal2 37766 5372 37766 5372 0 _0011_
rlabel metal2 42366 5032 42366 5032 0 _0012_
rlabel metal1 42964 3094 42964 3094 0 _0013_
rlabel via1 45030 4182 45030 4182 0 _0014_
rlabel metal1 39192 3094 39192 3094 0 _0015_
rlabel metal1 36984 4182 36984 4182 0 _0016_
rlabel metal1 35420 3094 35420 3094 0 _0017_
rlabel metal2 41262 4590 41262 4590 0 _0018_
rlabel metal2 40802 6698 40802 6698 0 _0019_
rlabel metal1 37398 3400 37398 3400 0 _0020_
rlabel metal1 22218 18938 22218 18938 0 _0021_
rlabel metal1 21804 18734 21804 18734 0 _0022_
rlabel metal1 46322 3570 46322 3570 0 _0023_
rlabel metal2 41998 23324 41998 23324 0 _0024_
rlabel metal2 53038 24004 53038 24004 0 _0025_
rlabel metal1 54970 22576 54970 22576 0 _0026_
rlabel metal2 55706 22746 55706 22746 0 _0027_
rlabel metal2 56534 16422 56534 16422 0 _0028_
rlabel metal2 56626 17238 56626 17238 0 _0029_
rlabel metal2 55614 22882 55614 22882 0 _0030_
rlabel metal2 56166 24276 56166 24276 0 _0031_
rlabel metal2 57086 25670 57086 25670 0 _0032_
rlabel metal1 58098 25840 58098 25840 0 _0033_
rlabel metal2 57914 26928 57914 26928 0 _0034_
rlabel metal1 57178 25976 57178 25976 0 _0035_
rlabel metal2 36386 6018 36386 6018 0 _0036_
rlabel metal2 55614 27812 55614 27812 0 _0037_
rlabel metal2 57224 25874 57224 25874 0 _0038_
rlabel metal2 56994 27914 56994 27914 0 _0039_
rlabel metal1 56442 22406 56442 22406 0 _0040_
rlabel metal1 52532 24106 52532 24106 0 _0041_
rlabel metal1 51198 17102 51198 17102 0 _0042_
rlabel metal2 53038 18768 53038 18768 0 _0043_
rlabel metal1 53268 20570 53268 20570 0 _0044_
rlabel metal1 55361 20910 55361 20910 0 _0045_
rlabel metal1 41124 2618 41124 2618 0 _0046_
rlabel metal2 53314 17136 53314 17136 0 _0047_
rlabel metal2 53130 19652 53130 19652 0 _0048_
rlabel metal1 55522 20434 55522 20434 0 _0049_
rlabel metal1 56718 20808 56718 20808 0 _0050_
rlabel metal1 56626 19346 56626 19346 0 _0051_
rlabel metal1 57040 21522 57040 21522 0 _0052_
rlabel metal2 56902 21318 56902 21318 0 _0053_
rlabel via1 56818 22678 56818 22678 0 _0054_
rlabel metal2 57454 22610 57454 22610 0 _0055_
rlabel metal2 56994 22882 56994 22882 0 _0056_
rlabel metal2 31786 14314 31786 14314 0 _0057_
rlabel metal1 57868 25330 57868 25330 0 _0058_
rlabel metal1 57822 25942 57822 25942 0 _0059_
rlabel metal1 57585 25262 57585 25262 0 _0060_
rlabel metal2 57546 20706 57546 20706 0 _0061_
rlabel metal2 51014 18326 51014 18326 0 _0062_
rlabel metal2 51106 19312 51106 19312 0 _0063_
rlabel metal1 56672 19278 56672 19278 0 _0064_
rlabel metal1 57316 19482 57316 19482 0 _0065_
rlabel metal1 57776 20026 57776 20026 0 _0066_
rlabel metal2 31786 7905 31786 7905 0 _0067_
rlabel metal2 58282 22583 58282 22583 0 _0068_
rlabel metal1 57868 24174 57868 24174 0 _0069_
rlabel metal2 58190 21828 58190 21828 0 _0070_
rlabel metal1 57132 23562 57132 23562 0 _0071_
rlabel metal1 57684 23494 57684 23494 0 _0072_
rlabel metal2 56350 24242 56350 24242 0 _0073_
rlabel metal1 56028 19754 56028 19754 0 _0074_
rlabel metal1 56488 23698 56488 23698 0 _0075_
rlabel metal2 56442 24004 56442 24004 0 _0076_
rlabel metal1 37720 6630 37720 6630 0 _0077_
rlabel metal1 58190 23290 58190 23290 0 _0078_
rlabel metal1 57224 24242 57224 24242 0 _0079_
rlabel metal2 56994 24378 56994 24378 0 _0080_
rlabel metal2 47702 4879 47702 4879 0 _0081_
rlabel metal2 40526 4250 40526 4250 0 _0082_
rlabel metal1 41538 6970 41538 6970 0 _0083_
rlabel metal1 32476 2550 32476 2550 0 _0084_
rlabel metal1 40848 3162 40848 3162 0 _0085_
rlabel metal2 41354 5236 41354 5236 0 _0086_
rlabel metal2 41446 7310 41446 7310 0 _0087_
rlabel metal1 41170 6800 41170 6800 0 _0088_
rlabel metal1 43524 7514 43524 7514 0 _0089_
rlabel metal1 35558 15028 35558 15028 0 _0090_
rlabel metal1 44850 5814 44850 5814 0 _0091_
rlabel metal1 45034 6698 45034 6698 0 _0092_
rlabel metal2 46322 6460 46322 6460 0 _0093_
rlabel metal1 40756 6426 40756 6426 0 _0094_
rlabel metal1 38548 5882 38548 5882 0 _0095_
rlabel metal1 41446 13872 41446 13872 0 _0096_
rlabel metal1 38824 5610 38824 5610 0 _0097_
rlabel metal2 40434 7888 40434 7888 0 _0098_
rlabel metal1 40250 9010 40250 9010 0 _0099_
rlabel metal1 22218 18700 22218 18700 0 _0100_
rlabel metal1 50692 4046 50692 4046 0 _0101_
rlabel metal1 47518 4114 47518 4114 0 _0102_
rlabel metal1 37766 15470 37766 15470 0 _0103_
rlabel metal1 42826 23664 42826 23664 0 _0104_
rlabel metal1 36938 16116 36938 16116 0 _0105_
rlabel metal2 31602 13401 31602 13401 0 _0106_
rlabel metal2 39238 14348 39238 14348 0 _0107_
rlabel metal1 32108 14586 32108 14586 0 _0108_
rlabel metal1 32223 12818 32223 12818 0 _0109_
rlabel metal2 32430 6902 32430 6902 0 _0110_
rlabel metal1 26818 13906 26818 13906 0 _0111_
rlabel metal1 32200 15470 32200 15470 0 _0112_
rlabel metal2 29946 15572 29946 15572 0 _0113_
rlabel via2 43654 19363 43654 19363 0 _0114_
rlabel metal1 43240 18734 43240 18734 0 _0115_
rlabel metal2 42826 19142 42826 19142 0 _0116_
rlabel metal2 27186 16218 27186 16218 0 _0117_
rlabel metal1 24380 14586 24380 14586 0 _0118_
rlabel metal1 23644 15130 23644 15130 0 _0119_
rlabel metal2 42642 20604 42642 20604 0 _0120_
rlabel metal2 22402 14858 22402 14858 0 _0121_
rlabel via2 28566 10421 28566 10421 0 _0122_
rlabel metal1 39054 12750 39054 12750 0 _0123_
rlabel metal1 24794 12818 24794 12818 0 _0124_
rlabel metal1 30176 6358 30176 6358 0 _0125_
rlabel metal1 31924 2822 31924 2822 0 _0126_
rlabel metal1 25530 9996 25530 9996 0 _0127_
rlabel metal1 30636 6358 30636 6358 0 _0128_
rlabel metal2 25346 5406 25346 5406 0 _0129_
rlabel metal2 39238 13600 39238 13600 0 _0130_
rlabel metal1 28750 5236 28750 5236 0 _0131_
rlabel metal1 30268 2550 30268 2550 0 _0132_
rlabel metal2 25990 8228 25990 8228 0 _0133_
rlabel metal1 29670 5236 29670 5236 0 _0134_
rlabel metal1 25438 12682 25438 12682 0 _0135_
rlabel metal1 36156 8466 36156 8466 0 _0136_
rlabel metal1 27876 6970 27876 6970 0 _0137_
rlabel metal1 28198 8976 28198 8976 0 _0138_
rlabel metal2 29578 5372 29578 5372 0 _0139_
rlabel metal3 29509 15300 29509 15300 0 _0140_
rlabel metal1 33902 8942 33902 8942 0 _0141_
rlabel metal2 33626 13124 33626 13124 0 _0142_
rlabel metal1 29164 12954 29164 12954 0 _0143_
rlabel metal2 32890 8466 32890 8466 0 _0144_
rlabel metal2 32154 8381 32154 8381 0 _0145_
rlabel metal1 32062 5100 32062 5100 0 _0146_
rlabel metal1 30084 15470 30084 15470 0 _0147_
rlabel metal1 28888 14994 28888 14994 0 _0148_
rlabel metal1 28888 15130 28888 15130 0 _0149_
rlabel metal2 28796 19210 28796 19210 0 _0150_
rlabel metal2 31648 23188 31648 23188 0 _0151_
rlabel metal1 38042 18632 38042 18632 0 _0152_
rlabel metal1 38640 13158 38640 13158 0 _0153_
rlabel metal1 29578 12818 29578 12818 0 _0154_
rlabel metal1 33994 2550 33994 2550 0 _0155_
rlabel metal1 34044 14382 34044 14382 0 _0156_
rlabel via2 28750 14059 28750 14059 0 _0157_
rlabel metal1 26174 13498 26174 13498 0 _0158_
rlabel metal1 28658 13328 28658 13328 0 _0159_
rlabel metal1 26726 12682 26726 12682 0 _0160_
rlabel metal1 26266 12852 26266 12852 0 _0161_
rlabel metal1 29900 13294 29900 13294 0 _0162_
rlabel metal1 29256 12614 29256 12614 0 _0163_
rlabel metal2 25898 13124 25898 13124 0 _0164_
rlabel metal1 25254 16966 25254 16966 0 _0165_
rlabel metal1 26358 22610 26358 22610 0 _0166_
rlabel metal1 35696 9146 35696 9146 0 _0167_
rlabel metal1 34040 7242 34040 7242 0 _0168_
rlabel metal2 32614 13328 32614 13328 0 _0169_
rlabel metal1 26496 5678 26496 5678 0 _0170_
rlabel metal1 32430 12410 32430 12410 0 _0171_
rlabel metal2 37122 5746 37122 5746 0 _0172_
rlabel metal1 33810 6766 33810 6766 0 _0173_
rlabel metal1 36202 12614 36202 12614 0 _0174_
rlabel metal1 27876 14994 27876 14994 0 _0175_
rlabel metal1 34270 9078 34270 9078 0 _0176_
rlabel metal2 36478 6613 36478 6613 0 _0177_
rlabel metal2 27462 7106 27462 7106 0 _0178_
rlabel metal2 31326 4454 31326 4454 0 _0179_
rlabel metal1 31004 6426 31004 6426 0 _0180_
rlabel metal1 37306 13906 37306 13906 0 _0181_
rlabel metal1 27278 14994 27278 14994 0 _0182_
rlabel metal2 26266 22814 26266 22814 0 _0183_
rlabel metal2 27094 23630 27094 23630 0 _0184_
rlabel metal2 27830 23868 27830 23868 0 _0185_
rlabel metal1 26358 20876 26358 20876 0 _0186_
rlabel metal1 31786 18700 31786 18700 0 _0187_
rlabel metal1 40986 13362 40986 13362 0 _0188_
rlabel metal2 26266 9486 26266 9486 0 _0189_
rlabel metal1 25806 8534 25806 8534 0 _0190_
rlabel metal1 37168 6834 37168 6834 0 _0191_
rlabel metal1 25852 11322 25852 11322 0 _0192_
rlabel metal2 28382 4386 28382 4386 0 _0193_
rlabel metal1 32936 3706 32936 3706 0 _0194_
rlabel via2 28014 4029 28014 4029 0 _0195_
rlabel metal1 27554 14450 27554 14450 0 _0196_
rlabel metal2 27462 11526 27462 11526 0 _0197_
rlabel metal1 24748 17170 24748 17170 0 _0198_
rlabel metal2 25622 18428 25622 18428 0 _0199_
rlabel metal2 26450 4386 26450 4386 0 _0200_
rlabel metal2 28934 7548 28934 7548 0 _0201_
rlabel metal2 27462 8228 27462 8228 0 _0202_
rlabel metal2 39422 10132 39422 10132 0 _0203_
rlabel metal1 27968 6698 27968 6698 0 _0204_
rlabel metal2 27370 5440 27370 5440 0 _0205_
rlabel metal1 38732 8262 38732 8262 0 _0206_
rlabel metal1 28060 5678 28060 5678 0 _0207_
rlabel metal1 27784 4794 27784 4794 0 _0208_
rlabel metal2 27186 7174 27186 7174 0 _0209_
rlabel metal1 26414 17578 26414 17578 0 _0210_
rlabel metal2 26358 18836 26358 18836 0 _0211_
rlabel metal2 26266 18836 26266 18836 0 _0212_
rlabel metal1 28842 11085 28842 11085 0 _0213_
rlabel metal1 28750 9588 28750 9588 0 _0214_
rlabel metal1 28704 8602 28704 8602 0 _0215_
rlabel metal1 40296 7378 40296 7378 0 _0216_
rlabel metal2 41078 8058 41078 8058 0 _0217_
rlabel metal1 28428 9622 28428 9622 0 _0218_
rlabel metal1 29670 9078 29670 9078 0 _0219_
rlabel metal1 27600 9622 27600 9622 0 _0220_
rlabel metal1 27186 9690 27186 9690 0 _0221_
rlabel metal2 26818 10336 26818 10336 0 _0222_
rlabel metal1 26818 15878 26818 15878 0 _0223_
rlabel metal1 26358 15674 26358 15674 0 _0224_
rlabel metal1 29072 16150 29072 16150 0 _0225_
rlabel via1 25425 7854 25425 7854 0 _0226_
rlabel metal2 24978 11526 24978 11526 0 _0227_
rlabel via2 33350 12291 33350 12291 0 _0228_
rlabel metal1 25116 14926 25116 14926 0 _0229_
rlabel metal2 25898 6324 25898 6324 0 _0230_
rlabel metal1 28152 6630 28152 6630 0 _0231_
rlabel via1 25162 6766 25162 6766 0 _0232_
rlabel metal1 25576 14994 25576 14994 0 _0233_
rlabel metal2 26450 15606 26450 15606 0 _0234_
rlabel metal1 29762 16558 29762 16558 0 _0235_
rlabel metal1 29946 16660 29946 16660 0 _0236_
rlabel metal1 27186 17170 27186 17170 0 _0237_
rlabel metal2 26266 16796 26266 16796 0 _0238_
rlabel metal2 26542 17986 26542 17986 0 _0239_
rlabel metal1 26174 20978 26174 20978 0 _0240_
rlabel metal2 37490 17918 37490 17918 0 _0241_
rlabel via1 26174 20893 26174 20893 0 _0242_
rlabel metal1 36386 18258 36386 18258 0 _0243_
rlabel metal1 36524 14314 36524 14314 0 _0244_
rlabel metal1 24978 8058 24978 8058 0 _0245_
rlabel metal1 34316 11118 34316 11118 0 _0246_
rlabel metal1 28290 9146 28290 9146 0 _0247_
rlabel metal2 25622 8670 25622 8670 0 _0248_
rlabel metal1 27646 19822 27646 19822 0 _0249_
rlabel metal1 29716 19346 29716 19346 0 _0250_
rlabel metal2 29762 20230 29762 20230 0 _0251_
rlabel metal1 37812 8942 37812 8942 0 _0252_
rlabel metal1 30452 7310 30452 7310 0 _0253_
rlabel metal2 30498 7548 30498 7548 0 _0254_
rlabel metal1 32614 6664 32614 6664 0 _0255_
rlabel metal1 30268 6834 30268 6834 0 _0256_
rlabel metal1 30314 7480 30314 7480 0 _0257_
rlabel metal1 38962 11118 38962 11118 0 _0258_
rlabel metal2 29302 11900 29302 11900 0 _0259_
rlabel metal1 29164 18734 29164 18734 0 _0260_
rlabel metal1 27094 20910 27094 20910 0 _0261_
rlabel metal2 24886 21760 24886 21760 0 _0262_
rlabel metal1 25392 21114 25392 21114 0 _0263_
rlabel metal2 24886 18020 24886 18020 0 _0264_
rlabel metal2 24794 17986 24794 17986 0 _0265_
rlabel metal2 25070 16830 25070 16830 0 _0266_
rlabel metal2 24058 18836 24058 18836 0 _0267_
rlabel metal2 25530 19686 25530 19686 0 _0268_
rlabel metal1 24012 20366 24012 20366 0 _0269_
rlabel metal2 23966 19210 23966 19210 0 _0270_
rlabel metal1 24242 21522 24242 21522 0 _0271_
rlabel metal2 23874 21386 23874 21386 0 _0272_
rlabel metal1 24656 21114 24656 21114 0 _0273_
rlabel metal2 23690 21318 23690 21318 0 _0274_
rlabel metal1 23552 20026 23552 20026 0 _0275_
rlabel metal1 23230 22542 23230 22542 0 _0276_
rlabel metal1 23598 23120 23598 23120 0 _0277_
rlabel metal2 23414 21726 23414 21726 0 _0278_
rlabel metal2 27094 21012 27094 21012 0 _0279_
rlabel metal2 27186 21828 27186 21828 0 _0280_
rlabel metal1 32798 17612 32798 17612 0 _0281_
rlabel metal1 28865 10778 28865 10778 0 _0282_
rlabel metal2 28290 11526 28290 11526 0 _0283_
rlabel metal2 28106 10234 28106 10234 0 _0284_
rlabel metal3 34017 9724 34017 9724 0 _0285_
rlabel metal2 33902 10370 33902 10370 0 _0286_
rlabel metal1 35926 13872 35926 13872 0 _0287_
rlabel metal1 28014 9996 28014 9996 0 _0288_
rlabel metal2 24794 10302 24794 10302 0 _0289_
rlabel metal2 24886 10234 24886 10234 0 _0290_
rlabel metal2 24702 10404 24702 10404 0 _0291_
rlabel metal1 27600 10030 27600 10030 0 _0292_
rlabel metal1 33074 18802 33074 18802 0 _0293_
rlabel metal1 28152 17510 28152 17510 0 _0294_
rlabel metal1 28152 17646 28152 17646 0 _0295_
rlabel metal2 26634 16388 26634 16388 0 _0296_
rlabel metal2 27738 12988 27738 12988 0 _0297_
rlabel metal2 27186 12308 27186 12308 0 _0298_
rlabel metal1 27324 12410 27324 12410 0 _0299_
rlabel metal1 28060 17170 28060 17170 0 _0300_
rlabel metal2 27646 16796 27646 16796 0 _0301_
rlabel metal2 28014 17170 28014 17170 0 _0302_
rlabel metal2 27922 19414 27922 19414 0 _0303_
rlabel via1 27838 20774 27838 20774 0 _0304_
rlabel metal1 28060 21114 28060 21114 0 _0305_
rlabel metal2 28106 19516 28106 19516 0 _0306_
rlabel metal2 33902 12002 33902 12002 0 _0307_
rlabel metal2 30084 13702 30084 13702 0 _0308_
rlabel metal2 29716 13124 29716 13124 0 _0309_
rlabel metal1 29440 11322 29440 11322 0 _0310_
rlabel metal1 28750 13260 28750 13260 0 _0311_
rlabel metal1 29302 13294 29302 13294 0 _0312_
rlabel metal2 30038 14518 30038 14518 0 _0313_
rlabel metal2 29670 16626 29670 16626 0 _0314_
rlabel metal1 27876 21454 27876 21454 0 _0315_
rlabel metal1 27692 21998 27692 21998 0 _0316_
rlabel metal1 28060 22542 28060 22542 0 _0317_
rlabel metal1 29854 23222 29854 23222 0 _0318_
rlabel metal1 28014 23290 28014 23290 0 _0319_
rlabel metal2 24518 21760 24518 21760 0 _0320_
rlabel metal1 29762 22610 29762 22610 0 _0321_
rlabel metal2 31602 19142 31602 19142 0 _0322_
rlabel metal1 33074 10064 33074 10064 0 _0323_
rlabel metal1 33396 9418 33396 9418 0 _0324_
rlabel metal1 33948 6970 33948 6970 0 _0325_
rlabel viali 33890 8466 33890 8466 0 _0326_
rlabel metal1 35006 8330 35006 8330 0 _0327_
rlabel metal1 33718 7854 33718 7854 0 _0328_
rlabel viali 32973 9554 32973 9554 0 _0329_
rlabel metal1 32660 17646 32660 17646 0 _0330_
rlabel metal2 31694 20230 31694 20230 0 _0331_
rlabel metal2 31786 19822 31786 19822 0 _0332_
rlabel metal2 31326 16252 31326 16252 0 _0333_
rlabel metal1 31050 15368 31050 15368 0 _0334_
rlabel metal1 32315 16082 32315 16082 0 _0335_
rlabel metal1 31096 16762 31096 16762 0 _0336_
rlabel metal1 31832 5338 31832 5338 0 _0337_
rlabel metal1 37122 16728 37122 16728 0 _0338_
rlabel metal1 30682 11118 30682 11118 0 _0339_
rlabel metal2 31786 10438 31786 10438 0 _0340_
rlabel metal1 31004 10778 31004 10778 0 _0341_
rlabel metal1 30958 9622 30958 9622 0 _0342_
rlabel metal1 30728 17170 30728 17170 0 _0343_
rlabel metal2 34178 16014 34178 16014 0 _0344_
rlabel metal2 31234 17510 31234 17510 0 _0345_
rlabel metal2 31418 19108 31418 19108 0 _0346_
rlabel metal2 31510 20842 31510 20842 0 _0347_
rlabel metal1 32292 20366 32292 20366 0 _0348_
rlabel viali 32798 6765 32798 6765 0 _0349_
rlabel metal2 32522 6681 32522 6681 0 _0350_
rlabel metal1 38548 12818 38548 12818 0 _0351_
rlabel metal2 35190 13022 35190 13022 0 _0352_
rlabel metal1 30820 9146 30820 9146 0 _0353_
rlabel metal2 31326 13770 31326 13770 0 _0354_
rlabel metal2 30406 16388 30406 16388 0 _0355_
rlabel metal1 29486 18938 29486 18938 0 _0356_
rlabel metal2 30038 18598 30038 18598 0 _0357_
rlabel metal1 30544 20434 30544 20434 0 _0358_
rlabel metal2 30682 21250 30682 21250 0 _0359_
rlabel metal1 30406 20910 30406 20910 0 _0360_
rlabel metal1 28290 20570 28290 20570 0 _0361_
rlabel metal1 30038 20876 30038 20876 0 _0362_
rlabel metal1 30222 22950 30222 22950 0 _0363_
rlabel metal1 30636 22610 30636 22610 0 _0364_
rlabel metal1 31418 23664 31418 23664 0 _0365_
rlabel metal2 29026 22916 29026 22916 0 _0366_
rlabel metal1 29992 23290 29992 23290 0 _0367_
rlabel metal1 57684 23698 57684 23698 0 _0368_
rlabel metal2 32338 21250 32338 21250 0 _0369_
rlabel metal1 35144 14994 35144 14994 0 _0370_
rlabel metal1 34040 14858 34040 14858 0 _0371_
rlabel metal1 32430 14042 32430 14042 0 _0372_
rlabel metal2 40434 9486 40434 9486 0 _0373_
rlabel metal1 32200 10778 32200 10778 0 _0374_
rlabel metal1 32246 11322 32246 11322 0 _0375_
rlabel metal2 32430 16116 32430 16116 0 _0376_
rlabel metal2 32522 19108 32522 19108 0 _0377_
rlabel metal1 33350 19754 33350 19754 0 _0378_
rlabel metal1 34132 14042 34132 14042 0 _0379_
rlabel metal1 33782 13906 33782 13906 0 _0380_
rlabel metal1 33304 15334 33304 15334 0 _0381_
rlabel metal1 33396 12954 33396 12954 0 _0382_
rlabel metal1 33120 13906 33120 13906 0 _0383_
rlabel metal1 33304 15470 33304 15470 0 _0384_
rlabel metal2 32798 15844 32798 15844 0 _0385_
rlabel metal1 33488 16218 33488 16218 0 _0386_
rlabel metal1 33120 16422 33120 16422 0 _0387_
rlabel metal1 34408 17714 34408 17714 0 _0388_
rlabel metal1 33718 19754 33718 19754 0 _0389_
rlabel via1 33718 21046 33718 21046 0 _0390_
rlabel metal1 33504 20842 33504 20842 0 _0391_
rlabel metal2 33350 21556 33350 21556 0 _0392_
rlabel metal1 35144 19822 35144 19822 0 _0393_
rlabel metal1 35374 20026 35374 20026 0 _0394_
rlabel metal1 38134 13362 38134 13362 0 _0395_
rlabel metal3 37260 9316 37260 9316 0 _0396_
rlabel metal2 36570 10676 36570 10676 0 _0397_
rlabel metal2 36662 6732 36662 6732 0 _0398_
rlabel metal1 36662 9690 36662 9690 0 _0399_
rlabel metal1 35788 20366 35788 20366 0 _0400_
rlabel metal1 34362 20910 34362 20910 0 _0401_
rlabel metal1 31786 21488 31786 21488 0 _0402_
rlabel metal2 30774 22644 30774 22644 0 _0403_
rlabel metal1 31372 23086 31372 23086 0 _0404_
rlabel metal2 32522 23664 32522 23664 0 _0405_
rlabel metal2 31602 24004 31602 24004 0 _0406_
rlabel metal1 38456 17578 38456 17578 0 _0407_
rlabel metal1 38456 17850 38456 17850 0 _0408_
rlabel metal1 40296 11050 40296 11050 0 _0409_
rlabel metal1 40250 11764 40250 11764 0 _0410_
rlabel metal2 40434 11322 40434 11322 0 _0411_
rlabel metal2 37582 9418 37582 9418 0 _0412_
rlabel metal1 37306 10574 37306 10574 0 _0413_
rlabel metal1 38594 10234 38594 10234 0 _0414_
rlabel metal1 40618 13158 40618 13158 0 _0415_
rlabel metal1 36524 13906 36524 13906 0 _0416_
rlabel metal1 40480 13362 40480 13362 0 _0417_
rlabel metal2 40342 15028 40342 15028 0 _0418_
rlabel metal1 40388 16762 40388 16762 0 _0419_
rlabel metal1 39744 16422 39744 16422 0 _0420_
rlabel metal2 36386 14722 36386 14722 0 _0421_
rlabel metal2 36202 8058 36202 8058 0 _0422_
rlabel metal1 35374 8058 35374 8058 0 _0423_
rlabel metal1 35742 8058 35742 8058 0 _0424_
rlabel metal1 35052 15402 35052 15402 0 _0425_
rlabel metal1 35098 15504 35098 15504 0 _0426_
rlabel metal2 35650 15844 35650 15844 0 _0427_
rlabel metal1 40526 16048 40526 16048 0 _0428_
rlabel metal1 40802 16218 40802 16218 0 _0429_
rlabel metal1 40572 17306 40572 17306 0 _0430_
rlabel metal2 41538 16320 41538 16320 0 _0431_
rlabel metal2 36754 18972 36754 18972 0 _0432_
rlabel metal2 36754 18496 36754 18496 0 _0433_
rlabel metal2 37766 11492 37766 11492 0 _0434_
rlabel metal1 37628 11866 37628 11866 0 _0435_
rlabel metal1 35420 13974 35420 13974 0 _0436_
rlabel metal2 37950 14790 37950 14790 0 _0437_
rlabel metal1 41814 16082 41814 16082 0 _0438_
rlabel metal1 36386 21964 36386 21964 0 _0439_
rlabel metal2 33810 21148 33810 21148 0 _0440_
rlabel metal2 35558 21760 35558 21760 0 _0441_
rlabel metal2 34822 22406 34822 22406 0 _0442_
rlabel metal2 32154 21828 32154 21828 0 _0443_
rlabel metal2 33994 22780 33994 22780 0 _0444_
rlabel metal1 38502 14382 38502 14382 0 _0445_
rlabel metal2 38962 8772 38962 8772 0 _0446_
rlabel metal1 39008 17170 39008 17170 0 _0447_
rlabel metal1 39330 18190 39330 18190 0 _0448_
rlabel metal1 39192 18258 39192 18258 0 _0449_
rlabel metal2 33442 12036 33442 12036 0 _0450_
rlabel metal1 33672 11866 33672 11866 0 _0451_
rlabel metal2 36754 10982 36754 10982 0 _0452_
rlabel metal1 34086 10540 34086 10540 0 _0453_
rlabel metal1 33810 10778 33810 10778 0 _0454_
rlabel metal1 33258 16626 33258 16626 0 _0455_
rlabel metal2 32798 17340 32798 17340 0 _0456_
rlabel metal2 33166 17782 33166 17782 0 _0457_
rlabel metal1 35903 18122 35903 18122 0 _0458_
rlabel metal1 39652 18938 39652 18938 0 _0459_
rlabel metal2 40158 19023 40158 19023 0 _0460_
rlabel metal1 40388 18802 40388 18802 0 _0461_
rlabel metal1 40158 12342 40158 12342 0 _0462_
rlabel metal1 39698 12682 39698 12682 0 _0463_
rlabel metal1 40526 14450 40526 14450 0 _0464_
rlabel metal2 40618 16660 40618 16660 0 _0465_
rlabel metal1 41262 18292 41262 18292 0 _0466_
rlabel metal2 41446 17238 41446 17238 0 _0467_
rlabel metal2 41170 18870 41170 18870 0 _0468_
rlabel metal2 41262 19958 41262 19958 0 _0469_
rlabel metal1 41078 22032 41078 22032 0 _0470_
rlabel metal2 41446 20060 41446 20060 0 _0471_
rlabel metal1 40526 21556 40526 21556 0 _0472_
rlabel metal2 40894 21794 40894 21794 0 _0473_
rlabel metal1 40710 22066 40710 22066 0 _0474_
rlabel metal1 41400 22406 41400 22406 0 _0475_
rlabel metal2 35328 10404 35328 10404 0 _0476_
rlabel metal1 37398 14042 37398 14042 0 _0477_
rlabel metal1 34730 11764 34730 11764 0 _0478_
rlabel metal1 35006 11322 35006 11322 0 _0479_
rlabel metal1 35144 11662 35144 11662 0 _0480_
rlabel metal1 35558 10710 35558 10710 0 _0481_
rlabel metal1 34868 10778 34868 10778 0 _0482_
rlabel metal1 35420 17306 35420 17306 0 _0483_
rlabel metal1 35282 19278 35282 19278 0 _0484_
rlabel metal1 36938 19346 36938 19346 0 _0485_
rlabel metal1 38180 16422 38180 16422 0 _0486_
rlabel metal1 36754 9010 36754 9010 0 _0487_
rlabel metal1 37398 9146 37398 9146 0 _0488_
rlabel metal1 37030 14994 37030 14994 0 _0489_
rlabel metal2 37398 15844 37398 15844 0 _0490_
rlabel metal1 36846 16694 36846 16694 0 _0491_
rlabel metal1 38226 18292 38226 18292 0 _0492_
rlabel metal2 38042 18870 38042 18870 0 _0493_
rlabel metal1 38502 20026 38502 20026 0 _0494_
rlabel metal2 36754 15844 36754 15844 0 _0495_
rlabel metal2 36846 17952 36846 17952 0 _0496_
rlabel metal1 36294 15504 36294 15504 0 _0497_
rlabel metal2 36938 19958 36938 19958 0 _0498_
rlabel metal2 36754 20060 36754 20060 0 _0499_
rlabel metal1 38778 19890 38778 19890 0 _0500_
rlabel metal1 39744 20434 39744 20434 0 _0501_
rlabel metal1 40296 19822 40296 19822 0 _0502_
rlabel metal2 41078 21012 41078 21012 0 _0503_
rlabel metal2 42182 21726 42182 21726 0 _0504_
rlabel metal2 39146 20672 39146 20672 0 _0505_
rlabel metal2 39054 21012 39054 21012 0 _0506_
rlabel metal1 36708 12410 36708 12410 0 _0507_
rlabel metal1 36340 12954 36340 12954 0 _0508_
rlabel metal1 36570 15130 36570 15130 0 _0509_
rlabel metal1 36202 15674 36202 15674 0 _0510_
rlabel metal1 35696 17306 35696 17306 0 _0511_
rlabel metal1 36524 20910 36524 20910 0 _0512_
rlabel metal1 38640 14042 38640 14042 0 _0513_
rlabel metal2 38410 15606 38410 15606 0 _0514_
rlabel metal2 37858 17544 37858 17544 0 _0515_
rlabel metal2 37582 19924 37582 19924 0 _0516_
rlabel metal1 38042 21488 38042 21488 0 _0517_
rlabel metal1 39008 15130 39008 15130 0 _0518_
rlabel metal1 38456 20910 38456 20910 0 _0519_
rlabel metal2 39330 21828 39330 21828 0 _0520_
rlabel metal1 40020 22066 40020 22066 0 _0521_
rlabel metal1 39882 22644 39882 22644 0 _0522_
rlabel metal2 40526 22916 40526 22916 0 _0523_
rlabel metal1 40526 20026 40526 20026 0 _0524_
rlabel metal1 41216 23698 41216 23698 0 _0525_
rlabel metal1 40388 21862 40388 21862 0 _0526_
rlabel metal2 40894 23290 40894 23290 0 _0527_
rlabel metal1 40526 23698 40526 23698 0 _0528_
rlabel metal1 37858 21114 37858 21114 0 _0529_
rlabel metal1 38456 21114 38456 21114 0 _0530_
rlabel metal1 34362 16422 34362 16422 0 _0531_
rlabel metal2 35558 20417 35558 20417 0 _0532_
rlabel metal1 37444 13498 37444 13498 0 _0533_
rlabel metal1 35696 14042 35696 14042 0 _0534_
rlabel metal2 35926 21318 35926 21318 0 _0535_
rlabel metal1 36708 21658 36708 21658 0 _0536_
rlabel metal1 37444 16966 37444 16966 0 _0537_
rlabel metal1 37398 17306 37398 17306 0 _0538_
rlabel metal1 36662 17850 36662 17850 0 _0539_
rlabel metal1 36984 23086 36984 23086 0 _0540_
rlabel metal1 35512 18394 35512 18394 0 _0541_
rlabel metal1 38410 23120 38410 23120 0 _0542_
rlabel metal1 38548 24174 38548 24174 0 _0543_
rlabel metal1 39100 23290 39100 23290 0 _0544_
rlabel metal1 40710 24208 40710 24208 0 _0545_
rlabel metal2 40066 25874 40066 25874 0 _0546_
rlabel metal2 39974 24310 39974 24310 0 _0547_
rlabel metal2 40250 25092 40250 25092 0 _0548_
rlabel metal1 40802 56814 40802 56814 0 _0549_
rlabel metal2 37490 24616 37490 24616 0 _0550_
rlabel metal1 37720 24582 37720 24582 0 _0551_
rlabel metal1 35512 14586 35512 14586 0 _0552_
rlabel metal1 34408 16218 34408 16218 0 _0553_
rlabel metal1 34822 19482 34822 19482 0 _0554_
rlabel metal2 35926 23494 35926 23494 0 _0555_
rlabel metal1 35788 23630 35788 23630 0 _0556_
rlabel metal2 36386 24276 36386 24276 0 _0557_
rlabel metal2 37214 25058 37214 25058 0 _0558_
rlabel metal2 38042 24718 38042 24718 0 _0559_
rlabel metal2 38226 25092 38226 25092 0 _0560_
rlabel metal1 38732 25330 38732 25330 0 _0561_
rlabel metal2 38962 26044 38962 26044 0 _0562_
rlabel metal1 35512 23494 35512 23494 0 _0563_
rlabel metal2 35282 24004 35282 24004 0 _0564_
rlabel metal1 37444 24038 37444 24038 0 _0565_
rlabel metal2 38410 24582 38410 24582 0 _0566_
rlabel metal1 39192 24650 39192 24650 0 _0567_
rlabel metal1 36248 24582 36248 24582 0 _0568_
rlabel metal1 51290 6222 51290 6222 0 _0569_
rlabel metal1 43332 13906 43332 13906 0 _0570_
rlabel metal2 53038 8228 53038 8228 0 _0571_
rlabel metal1 42320 11662 42320 11662 0 _0572_
rlabel metal1 43240 12818 43240 12818 0 _0573_
rlabel metal2 45862 4964 45862 4964 0 _0574_
rlabel metal1 42136 8466 42136 8466 0 _0575_
rlabel metal1 41584 8330 41584 8330 0 _0576_
rlabel metal1 47794 13260 47794 13260 0 _0577_
rlabel metal2 47426 15810 47426 15810 0 _0578_
rlabel metal1 44574 16048 44574 16048 0 _0579_
rlabel metal1 48024 13294 48024 13294 0 _0580_
rlabel metal1 44804 16150 44804 16150 0 _0581_
rlabel metal2 44758 16388 44758 16388 0 _0582_
rlabel metal1 46046 8840 46046 8840 0 _0583_
rlabel metal2 46874 13974 46874 13974 0 _0584_
rlabel metal2 50462 13668 50462 13668 0 _0585_
rlabel metal1 46690 10234 46690 10234 0 _0586_
rlabel metal1 43240 13974 43240 13974 0 _0587_
rlabel metal1 53958 9962 53958 9962 0 _0588_
rlabel metal1 52118 8840 52118 8840 0 _0589_
rlabel metal1 56580 6834 56580 6834 0 _0590_
rlabel metal1 55384 6834 55384 6834 0 _0591_
rlabel metal1 51474 10472 51474 10472 0 _0592_
rlabel metal1 46966 10710 46966 10710 0 _0593_
rlabel metal2 46506 13532 46506 13532 0 _0594_
rlabel metal2 56810 16082 56810 16082 0 _0595_
rlabel metal1 44850 21862 44850 21862 0 _0596_
rlabel metal2 44482 23596 44482 23596 0 _0597_
rlabel metal2 58098 11866 58098 11866 0 _0598_
rlabel metal1 49450 13226 49450 13226 0 _0599_
rlabel metal1 53820 5270 53820 5270 0 _0600_
rlabel metal1 49634 17680 49634 17680 0 _0601_
rlabel via1 45769 16082 45769 16082 0 _0602_
rlabel metal2 47978 14484 47978 14484 0 _0603_
rlabel metal1 48668 13906 48668 13906 0 _0604_
rlabel metal1 46736 15470 46736 15470 0 _0605_
rlabel metal1 46000 15674 46000 15674 0 _0606_
rlabel metal1 43378 14382 43378 14382 0 _0607_
rlabel metal1 44413 13294 44413 13294 0 _0608_
rlabel metal1 42826 14586 42826 14586 0 _0609_
rlabel metal1 48346 13192 48346 13192 0 _0610_
rlabel metal1 44850 17136 44850 17136 0 _0611_
rlabel via2 44942 15011 44942 15011 0 _0612_
rlabel metal2 51106 7514 51106 7514 0 _0613_
rlabel metal1 51244 15062 51244 15062 0 _0614_
rlabel metal2 44666 16150 44666 16150 0 _0615_
rlabel metal2 45586 16558 45586 16558 0 _0616_
rlabel metal1 46000 22610 46000 22610 0 _0617_
rlabel via1 44290 26282 44290 26282 0 _0618_
rlabel metal1 47978 17850 47978 17850 0 _0619_
rlabel metal1 46092 8466 46092 8466 0 _0620_
rlabel metal1 48576 17850 48576 17850 0 _0621_
rlabel metal1 51244 16150 51244 16150 0 _0622_
rlabel metal2 52946 13260 52946 13260 0 _0623_
rlabel metal1 48254 18054 48254 18054 0 _0624_
rlabel metal2 47610 18428 47610 18428 0 _0625_
rlabel viali 47150 8471 47150 8471 0 _0626_
rlabel metal1 54372 8942 54372 8942 0 _0627_
rlabel metal2 47150 15844 47150 15844 0 _0628_
rlabel metal1 52256 4522 52256 4522 0 _0629_
rlabel metal2 58098 14144 58098 14144 0 _0630_
rlabel metal1 53958 9554 53958 9554 0 _0631_
rlabel metal2 47058 14586 47058 14586 0 _0632_
rlabel metal2 52118 9350 52118 9350 0 _0633_
rlabel metal1 47334 14042 47334 14042 0 _0634_
rlabel metal1 47702 14382 47702 14382 0 _0635_
rlabel metal2 46966 16660 46966 16660 0 _0636_
rlabel metal1 46276 19890 46276 19890 0 _0637_
rlabel metal1 43976 26826 43976 26826 0 _0638_
rlabel metal2 43838 24480 43838 24480 0 _0639_
rlabel metal1 52900 25806 52900 25806 0 _0640_
rlabel metal1 44068 26962 44068 26962 0 _0641_
rlabel metal2 44666 27778 44666 27778 0 _0642_
rlabel metal1 54142 21556 54142 21556 0 _0643_
rlabel metal1 48254 12172 48254 12172 0 _0644_
rlabel metal1 50186 6222 50186 6222 0 _0645_
rlabel metal2 55430 10472 55430 10472 0 _0646_
rlabel metal1 48852 8330 48852 8330 0 _0647_
rlabel metal1 47012 8602 47012 8602 0 _0648_
rlabel metal2 46230 9010 46230 9010 0 _0649_
rlabel metal1 51796 12750 51796 12750 0 _0650_
rlabel metal2 51566 10642 51566 10642 0 _0651_
rlabel metal2 46322 8993 46322 8993 0 _0652_
rlabel metal2 46644 17204 46644 17204 0 _0653_
rlabel metal1 46000 26554 46000 26554 0 _0654_
rlabel metal1 54188 9418 54188 9418 0 _0655_
rlabel metal1 46230 18326 46230 18326 0 _0656_
rlabel metal1 50324 9962 50324 9962 0 _0657_
rlabel metal2 48714 9860 48714 9860 0 _0658_
rlabel metal2 49910 6596 49910 6596 0 _0659_
rlabel metal2 54878 13396 54878 13396 0 _0660_
rlabel metal1 49496 6970 49496 6970 0 _0661_
rlabel metal1 52348 13906 52348 13906 0 _0662_
rlabel metal1 51934 14994 51934 14994 0 _0663_
rlabel metal1 49266 6800 49266 6800 0 _0664_
rlabel metal2 53406 7089 53406 7089 0 _0665_
rlabel metal2 49358 7004 49358 7004 0 _0666_
rlabel metal2 49082 8432 49082 8432 0 _0667_
rlabel metal2 48162 12342 48162 12342 0 _0668_
rlabel metal1 47472 22406 47472 22406 0 _0669_
rlabel metal2 45862 27744 45862 27744 0 _0670_
rlabel metal2 45770 27778 45770 27778 0 _0671_
rlabel metal1 46782 12614 46782 12614 0 _0672_
rlabel metal1 51842 16762 51842 16762 0 _0673_
rlabel metal1 47978 7820 47978 7820 0 _0674_
rlabel metal1 43240 11322 43240 11322 0 _0675_
rlabel metal1 44666 11798 44666 11798 0 _0676_
rlabel metal1 45632 14042 45632 14042 0 _0677_
rlabel metal1 45770 11662 45770 11662 0 _0678_
rlabel metal2 46874 12002 46874 12002 0 _0679_
rlabel metal1 46368 11186 46368 11186 0 _0680_
rlabel metal2 48070 10846 48070 10846 0 _0681_
rlabel metal2 47058 11356 47058 11356 0 _0682_
rlabel metal1 46230 19278 46230 19278 0 _0683_
rlabel metal1 48530 20366 48530 20366 0 _0684_
rlabel metal1 47058 20026 47058 20026 0 _0685_
rlabel metal1 49588 12886 49588 12886 0 _0686_
rlabel metal1 50692 13294 50692 13294 0 _0687_
rlabel metal1 50278 13226 50278 13226 0 _0688_
rlabel metal2 53866 13668 53866 13668 0 _0689_
rlabel via1 49266 12799 49266 12799 0 _0690_
rlabel metal2 49634 12410 49634 12410 0 _0691_
rlabel metal1 49082 19414 49082 19414 0 _0692_
rlabel metal2 44390 20196 44390 20196 0 _0693_
rlabel metal1 45356 20434 45356 20434 0 _0694_
rlabel metal1 45816 19754 45816 19754 0 _0695_
rlabel metal2 47794 21862 47794 21862 0 _0696_
rlabel metal1 46230 27438 46230 27438 0 _0697_
rlabel metal1 46391 28662 46391 28662 0 _0698_
rlabel metal2 46874 28764 46874 28764 0 _0699_
rlabel metal2 58006 6494 58006 6494 0 _0700_
rlabel metal1 44942 11866 44942 11866 0 _0701_
rlabel metal2 56718 8704 56718 8704 0 _0702_
rlabel metal2 44942 12036 44942 12036 0 _0703_
rlabel metal3 43999 18020 43999 18020 0 _0704_
rlabel metal1 43194 15436 43194 15436 0 _0705_
rlabel metal1 44390 17646 44390 17646 0 _0706_
rlabel metal1 44896 17850 44896 17850 0 _0707_
rlabel metal1 44206 18394 44206 18394 0 _0708_
rlabel metal1 45126 9622 45126 9622 0 _0709_
rlabel metal1 44666 7514 44666 7514 0 _0710_
rlabel metal2 44022 9078 44022 9078 0 _0711_
rlabel metal1 44100 9350 44100 9350 0 _0712_
rlabel metal1 43608 10030 43608 10030 0 _0713_
rlabel metal1 43516 10234 43516 10234 0 _0714_
rlabel metal3 43884 9724 43884 9724 0 _0715_
rlabel metal2 44896 18836 44896 18836 0 _0716_
rlabel metal1 44436 22202 44436 22202 0 _0717_
rlabel metal1 45908 28458 45908 28458 0 _0718_
rlabel metal1 47012 29138 47012 29138 0 _0719_
rlabel metal1 46184 28934 46184 28934 0 _0720_
rlabel metal1 45586 24786 45586 24786 0 _0721_
rlabel metal2 45586 23970 45586 23970 0 _0722_
rlabel metal1 46276 18938 46276 18938 0 _0723_
rlabel metal1 45816 19142 45816 19142 0 _0724_
rlabel metal1 45356 25466 45356 25466 0 _0725_
rlabel via1 45394 24106 45394 24106 0 _0726_
rlabel metal1 44758 29138 44758 29138 0 _0727_
rlabel metal2 43930 25636 43930 25636 0 _0728_
rlabel metal2 44758 27540 44758 27540 0 _0729_
rlabel metal1 46598 29648 46598 29648 0 _0730_
rlabel metal2 46782 30566 46782 30566 0 _0731_
rlabel via1 46414 29750 46414 29750 0 _0732_
rlabel metal1 47196 29818 47196 29818 0 _0733_
rlabel metal2 46966 30906 46966 30906 0 _0734_
rlabel metal2 44850 30804 44850 30804 0 _0735_
rlabel metal1 45034 30090 45034 30090 0 _0736_
rlabel metal1 46230 30294 46230 30294 0 _0737_
rlabel metal1 46828 25874 46828 25874 0 _0738_
rlabel metal2 46322 7582 46322 7582 0 _0739_
rlabel metal1 46506 5882 46506 5882 0 _0740_
rlabel metal1 46897 7378 46897 7378 0 _0741_
rlabel metal1 47242 7310 47242 7310 0 _0742_
rlabel metal1 45908 7514 45908 7514 0 _0743_
rlabel metal1 42182 10132 42182 10132 0 _0744_
rlabel metal1 45310 10132 45310 10132 0 _0745_
rlabel via2 45954 10251 45954 10251 0 _0746_
rlabel metal2 48070 26146 48070 26146 0 _0747_
rlabel metal1 48162 26418 48162 26418 0 _0748_
rlabel metal1 48484 20910 48484 20910 0 _0749_
rlabel metal1 46322 20434 46322 20434 0 _0750_
rlabel metal1 51888 20910 51888 20910 0 _0751_
rlabel metal2 42734 14518 42734 14518 0 _0752_
rlabel metal1 44252 15878 44252 15878 0 _0753_
rlabel metal1 47940 15130 47940 15130 0 _0754_
rlabel metal2 48530 15487 48530 15487 0 _0755_
rlabel metal2 48530 16320 48530 16320 0 _0756_
rlabel metal1 48208 20434 48208 20434 0 _0757_
rlabel metal1 47656 20978 47656 20978 0 _0758_
rlabel metal2 47518 21563 47518 21563 0 _0759_
rlabel metal1 47518 26554 47518 26554 0 _0760_
rlabel metal1 48162 27098 48162 27098 0 _0761_
rlabel metal1 47886 27506 47886 27506 0 _0762_
rlabel metal1 45908 6766 45908 6766 0 _0763_
rlabel metal1 52624 9418 52624 9418 0 _0764_
rlabel metal2 51934 11220 51934 11220 0 _0765_
rlabel metal2 53866 16354 53866 16354 0 _0766_
rlabel metal2 50830 11968 50830 11968 0 _0767_
rlabel metal2 51658 10438 51658 10438 0 _0768_
rlabel metal1 51520 11730 51520 11730 0 _0769_
rlabel metal2 50646 12342 50646 12342 0 _0770_
rlabel metal1 50232 12954 50232 12954 0 _0771_
rlabel metal1 48162 24718 48162 24718 0 _0772_
rlabel metal1 47564 24922 47564 24922 0 _0773_
rlabel metal1 47656 27506 47656 27506 0 _0774_
rlabel metal2 47978 28356 47978 28356 0 _0775_
rlabel metal2 48162 29342 48162 29342 0 _0776_
rlabel metal2 49266 29954 49266 29954 0 _0777_
rlabel metal1 49266 28560 49266 28560 0 _0778_
rlabel metal1 48622 29818 48622 29818 0 _0779_
rlabel metal2 48346 30498 48346 30498 0 _0780_
rlabel metal2 52210 23392 52210 23392 0 _0781_
rlabel metal2 46782 23188 46782 23188 0 _0782_
rlabel metal2 50186 14178 50186 14178 0 _0783_
rlabel metal2 41446 14824 41446 14824 0 _0784_
rlabel metal2 45724 14586 45724 14586 0 _0785_
rlabel metal1 42964 14518 42964 14518 0 _0786_
rlabel metal2 45678 15164 45678 15164 0 _0787_
rlabel metal1 45402 14926 45402 14926 0 _0788_
rlabel metal2 48714 23290 48714 23290 0 _0789_
rlabel metal1 48944 20910 48944 20910 0 _0790_
rlabel metal1 53176 10234 53176 10234 0 _0791_
rlabel metal1 54004 10234 54004 10234 0 _0792_
rlabel metal1 55844 11322 55844 11322 0 _0793_
rlabel metal1 55016 11186 55016 11186 0 _0794_
rlabel via2 51382 16541 51382 16541 0 _0795_
rlabel metal1 51658 16218 51658 16218 0 _0796_
rlabel metal1 50968 11322 50968 11322 0 _0797_
rlabel metal1 51750 16490 51750 16490 0 _0798_
rlabel via2 49174 20893 49174 20893 0 _0799_
rlabel metal1 49036 21114 49036 21114 0 _0800_
rlabel metal2 48806 21828 48806 21828 0 _0801_
rlabel metal1 49220 10506 49220 10506 0 _0802_
rlabel metal2 54234 13668 54234 13668 0 _0803_
rlabel metal1 48392 8058 48392 8058 0 _0804_
rlabel metal1 48438 11866 48438 11866 0 _0805_
rlabel metal2 49450 11798 49450 11798 0 _0806_
rlabel metal1 48530 11322 48530 11322 0 _0807_
rlabel metal1 49036 19210 49036 19210 0 _0808_
rlabel metal1 51704 20978 51704 20978 0 _0809_
rlabel metal1 49404 22066 49404 22066 0 _0810_
rlabel metal2 48990 23426 48990 23426 0 _0811_
rlabel metal2 49174 24480 49174 24480 0 _0812_
rlabel metal2 49266 24650 49266 24650 0 _0813_
rlabel metal1 54004 13838 54004 13838 0 _0814_
rlabel viali 48988 14994 48988 14994 0 _0815_
rlabel metal2 48898 14756 48898 14756 0 _0816_
rlabel metal1 51980 20230 51980 20230 0 _0817_
rlabel metal1 48806 14382 48806 14382 0 _0818_
rlabel metal1 43608 14042 43608 14042 0 _0819_
rlabel metal1 48116 14382 48116 14382 0 _0820_
rlabel metal2 48070 14790 48070 14790 0 _0821_
rlabel metal2 48530 25041 48530 25041 0 _0822_
rlabel metal1 48990 25330 48990 25330 0 _0823_
rlabel metal1 49404 25942 49404 25942 0 _0824_
rlabel metal1 45034 13906 45034 13906 0 _0825_
rlabel metal1 49588 27302 49588 27302 0 _0826_
rlabel metal2 49726 26996 49726 26996 0 _0827_
rlabel metal1 49358 28016 49358 28016 0 _0828_
rlabel metal1 51796 28526 51796 28526 0 _0829_
rlabel metal2 49634 28900 49634 28900 0 _0830_
rlabel metal1 51566 28560 51566 28560 0 _0831_
rlabel metal2 49450 29274 49450 29274 0 _0832_
rlabel metal1 50186 28526 50186 28526 0 _0833_
rlabel via2 47058 2635 47058 2635 0 _0834_
rlabel metal2 54602 14144 54602 14144 0 _0835_
rlabel metal1 50324 27030 50324 27030 0 _0836_
rlabel metal2 46690 23494 46690 23494 0 _0837_
rlabel metal1 45540 17714 45540 17714 0 _0838_
rlabel metal1 46138 12954 46138 12954 0 _0839_
rlabel metal2 46414 15079 46414 15079 0 _0840_
rlabel metal2 49818 17884 49818 17884 0 _0841_
rlabel metal1 49358 17510 49358 17510 0 _0842_
rlabel metal1 46598 17306 46598 17306 0 _0843_
rlabel metal2 46966 23902 46966 23902 0 _0844_
rlabel metal1 47564 23494 47564 23494 0 _0845_
rlabel metal2 54694 15300 54694 15300 0 _0846_
rlabel metal1 47434 23834 47434 23834 0 _0847_
rlabel metal1 49726 23766 49726 23766 0 _0848_
rlabel metal2 49174 20128 49174 20128 0 _0849_
rlabel metal1 49588 20502 49588 20502 0 _0850_
rlabel metal1 50002 23290 50002 23290 0 _0851_
rlabel metal1 50048 24786 50048 24786 0 _0852_
rlabel metal1 50784 25262 50784 25262 0 _0853_
rlabel metal1 51290 23732 51290 23732 0 _0854_
rlabel metal2 50830 24004 50830 24004 0 _0855_
rlabel metal1 52762 15470 52762 15470 0 _0856_
rlabel metal2 56166 9860 56166 9860 0 _0857_
rlabel metal1 52624 15062 52624 15062 0 _0858_
rlabel metal1 52348 14858 52348 14858 0 _0859_
rlabel metal2 47886 6256 47886 6256 0 _0860_
rlabel metal1 50646 14008 50646 14008 0 _0861_
rlabel metal1 53498 14416 53498 14416 0 _0862_
rlabel metal1 52992 14586 52992 14586 0 _0863_
rlabel metal1 51566 23698 51566 23698 0 _0864_
rlabel metal1 50692 25330 50692 25330 0 _0865_
rlabel metal1 50876 26282 50876 26282 0 _0866_
rlabel metal2 50922 28509 50922 28509 0 _0867_
rlabel metal1 56994 20230 56994 20230 0 _0868_
rlabel metal2 51152 27982 51152 27982 0 _0869_
rlabel metal2 51842 29444 51842 29444 0 _0870_
rlabel metal1 51244 29682 51244 29682 0 _0871_
rlabel metal2 51382 28288 51382 28288 0 _0872_
rlabel metal1 55844 12070 55844 12070 0 _0873_
rlabel metal1 55798 12206 55798 12206 0 _0874_
rlabel metal2 55982 12070 55982 12070 0 _0875_
rlabel metal3 53521 16660 53521 16660 0 _0876_
rlabel metal1 46506 18190 46506 18190 0 _0877_
rlabel metal1 55108 8466 55108 8466 0 _0878_
rlabel metal1 51796 17850 51796 17850 0 _0879_
rlabel metal1 53360 19278 53360 19278 0 _0880_
rlabel metal2 52118 22916 52118 22916 0 _0881_
rlabel metal1 45586 18122 45586 18122 0 _0882_
rlabel metal2 43470 16150 43470 16150 0 _0883_
rlabel metal1 43240 17306 43240 17306 0 _0884_
rlabel metal1 43700 17306 43700 17306 0 _0885_
rlabel metal1 44390 17782 44390 17782 0 _0886_
rlabel metal2 46414 18564 46414 18564 0 _0887_
rlabel metal1 52080 22950 52080 22950 0 _0888_
rlabel metal1 55936 9622 55936 9622 0 _0889_
rlabel metal1 52440 24786 52440 24786 0 _0890_
rlabel metal2 53222 24038 53222 24038 0 _0891_
rlabel metal1 53130 25262 53130 25262 0 _0892_
rlabel metal1 51796 23494 51796 23494 0 _0893_
rlabel metal1 53682 18700 53682 18700 0 _0894_
rlabel metal1 51520 14450 51520 14450 0 _0895_
rlabel metal1 51658 14042 51658 14042 0 _0896_
rlabel metal2 52578 15215 52578 15215 0 _0897_
rlabel metal2 52854 25058 52854 25058 0 _0898_
rlabel metal1 52302 25330 52302 25330 0 _0899_
rlabel metal1 54234 7174 54234 7174 0 _0900_
rlabel metal2 52210 26013 52210 26013 0 _0901_
rlabel metal2 52946 28016 52946 28016 0 _0902_
rlabel metal1 53176 28050 53176 28050 0 _0903_
rlabel metal1 51888 28050 51888 28050 0 _0904_
rlabel metal2 53222 27336 53222 27336 0 _0905_
rlabel metal2 53406 26656 53406 26656 0 _0906_
rlabel metal1 54234 12410 54234 12410 0 _0907_
rlabel metal2 53406 19516 53406 19516 0 _0908_
rlabel metal2 54418 14790 54418 14790 0 _0909_
rlabel metal1 55016 13158 55016 13158 0 _0910_
rlabel metal1 54372 21998 54372 21998 0 _0911_
rlabel metal1 54004 22066 54004 22066 0 _0912_
rlabel metal1 52992 21998 52992 21998 0 _0913_
rlabel metal1 50140 15334 50140 15334 0 _0914_
rlabel metal1 50738 15674 50738 15674 0 _0915_
rlabel metal1 52118 10778 52118 10778 0 _0916_
rlabel metal1 52164 11186 52164 11186 0 _0917_
rlabel metal2 54602 11186 54602 11186 0 _0918_
rlabel via1 51106 11237 51106 11237 0 _0919_
rlabel metal1 50094 16218 50094 16218 0 _0920_
rlabel metal1 54142 6324 54142 6324 0 _0921_
rlabel metal2 50186 21250 50186 21250 0 _0922_
rlabel metal1 53820 22610 53820 22610 0 _0923_
rlabel metal1 53452 23290 53452 23290 0 _0924_
rlabel metal1 54142 22644 54142 22644 0 _0925_
rlabel metal1 53820 23290 53820 23290 0 _0926_
rlabel metal1 53452 8942 53452 8942 0 _0927_
rlabel metal1 53728 9146 53728 9146 0 _0928_
rlabel via3 54027 18020 54027 18020 0 _0929_
rlabel metal1 54096 24174 54096 24174 0 _0930_
rlabel metal1 54188 25262 54188 25262 0 _0931_
rlabel metal1 46184 8058 46184 8058 0 _0932_
rlabel metal1 53038 24752 53038 24752 0 _0933_
rlabel metal1 53958 25296 53958 25296 0 _0934_
rlabel metal1 54050 25840 54050 25840 0 _0935_
rlabel metal1 54280 25874 54280 25874 0 _0936_
rlabel metal2 54050 26180 54050 26180 0 _0937_
rlabel metal1 52900 27098 52900 27098 0 _0938_
rlabel metal2 53958 27370 53958 27370 0 _0939_
rlabel metal2 53866 27370 53866 27370 0 _0940_
rlabel metal1 52716 12614 52716 12614 0 _0941_
rlabel metal1 46230 16490 46230 16490 0 _0942_
rlabel metal1 53498 12614 53498 12614 0 _0943_
rlabel metal1 53268 12410 53268 12410 0 _0944_
rlabel metal2 51382 10234 51382 10234 0 _0945_
rlabel metal1 52854 9962 52854 9962 0 _0946_
rlabel via2 52026 19261 52026 19261 0 _0947_
rlabel metal2 51382 20196 51382 20196 0 _0948_
rlabel metal1 51474 20400 51474 20400 0 _0949_
rlabel metal2 55522 24480 55522 24480 0 _0950_
rlabel metal1 52486 16626 52486 16626 0 _0951_
rlabel metal1 53176 16762 53176 16762 0 _0952_
rlabel metal2 55522 14484 55522 14484 0 _0953_
rlabel metal1 53590 17646 53590 17646 0 _0954_
rlabel metal2 54510 18836 54510 18836 0 _0955_
rlabel metal1 54372 20026 54372 20026 0 _0956_
rlabel metal1 55706 24140 55706 24140 0 _0957_
rlabel metal2 56442 25469 56442 25469 0 _0958_
rlabel metal1 53590 18224 53590 18224 0 _0959_
rlabel metal2 55154 18564 55154 18564 0 _0960_
rlabel metal1 56120 18598 56120 18598 0 _0961_
rlabel metal2 55522 19108 55522 19108 0 _0962_
rlabel metal2 56534 26418 56534 26418 0 _0963_
rlabel metal2 56074 27506 56074 27506 0 _0964_
rlabel metal2 53130 24004 53130 24004 0 _0965_
rlabel metal2 55890 27506 55890 27506 0 _0966_
rlabel metal2 55246 28560 55246 28560 0 _0967_
rlabel metal2 54418 27574 54418 27574 0 _0968_
rlabel metal2 54142 28288 54142 28288 0 _0969_
rlabel metal2 55890 25534 55890 25534 0 _0970_
rlabel metal1 55660 25670 55660 25670 0 _0971_
rlabel metal1 53498 14042 53498 14042 0 _0972_
rlabel metal1 39422 7922 39422 7922 0 _0973_
rlabel metal2 53774 17544 53774 17544 0 _0974_
rlabel metal2 53958 17782 53958 17782 0 _0975_
rlabel metal1 53130 18394 53130 18394 0 _0976_
rlabel metal1 51428 20026 51428 20026 0 _0977_
rlabel metal2 55246 21046 55246 21046 0 _0978_
rlabel metal2 54878 16966 54878 16966 0 _0979_
rlabel metal1 54510 20910 54510 20910 0 _0980_
rlabel metal1 54280 21114 54280 21114 0 _0981_
rlabel metal2 55062 21726 55062 21726 0 _0982_
rlabel metal1 55890 21862 55890 21862 0 _0983_
rlabel metal2 38318 6732 38318 6732 0 _0984_
rlabel metal2 16790 1520 16790 1520 0 addI[0]
rlabel metal2 21942 1520 21942 1520 0 addI[1]
rlabel metal2 58282 18513 58282 18513 0 addI[2]
rlabel metal2 27738 1520 27738 1520 0 addI[3]
rlabel via2 58282 54485 58282 54485 0 addI[4]
rlabel metal2 58282 58735 58282 58735 0 addI[5]
rlabel metal1 21712 57562 21712 57562 0 addQ[0]
rlabel metal1 26864 57562 26864 57562 0 addQ[1]
rlabel metal2 38686 1520 38686 1520 0 addQ[2]
rlabel metal3 1188 23188 1188 23188 0 addQ[3]
rlabel metal1 2254 57562 2254 57562 0 addQ[4]
rlabel via2 58282 24565 58282 24565 0 addQ[5]
rlabel metal2 48024 4522 48024 4522 0 bit2symb.regi
rlabel metal1 40940 2346 40940 2346 0 clknet_0_CLK
rlabel metal2 37490 2621 37490 2621 0 clknet_1_0__leaf_CLK
rlabel metal1 43562 2618 43562 2618 0 clknet_1_1__leaf_CLK
rlabel metal2 1794 11645 1794 11645 0 net1
rlabel metal1 49358 56678 49358 56678 0 net10
rlabel metal1 36294 2482 36294 2482 0 net11
rlabel metal1 57822 42670 57822 42670 0 net12
rlabel metal2 58098 7174 58098 7174 0 net13
rlabel metal1 12236 2414 12236 2414 0 net14
rlabel metal1 2116 41106 2116 41106 0 net15
rlabel metal2 2438 28424 2438 28424 0 net16
rlabel metal1 38134 57460 38134 57460 0 net17
rlabel metal1 41354 56712 41354 56712 0 net18
rlabel metal1 1932 35666 1932 35666 0 net19
rlabel metal1 32292 57358 32292 57358 0 net2
rlabel metal1 57178 25432 57178 25432 0 net20
rlabel metal1 19366 22950 19366 22950 0 net21
rlabel metal1 2162 2414 2162 2414 0 net22
rlabel metal1 24518 23630 24518 23630 0 net23
rlabel metal1 58144 30702 58144 30702 0 net24
rlabel metal1 10304 57426 10304 57426 0 net25
rlabel metal1 2162 5678 2162 5678 0 net26
rlabel metal1 50646 2448 50646 2448 0 net27
rlabel metal1 43884 57222 43884 57222 0 net28
rlabel metal1 58052 13294 58052 13294 0 net29
rlabel metal2 21390 14892 21390 14892 0 net3
rlabel metal2 17710 2176 17710 2176 0 net30
rlabel metal1 52072 2618 52072 2618 0 net31
rlabel metal1 58236 18734 58236 18734 0 net32
rlabel metal1 54832 13430 54832 13430 0 net33
rlabel metal1 57454 54502 57454 54502 0 net34
rlabel metal1 57638 57222 57638 57222 0 net35
rlabel metal1 22724 57222 22724 57222 0 net36
rlabel via2 28014 57205 28014 57205 0 net37
rlabel metal1 35190 3434 35190 3434 0 net38
rlabel metal1 2116 23698 2116 23698 0 net39
rlabel metal1 2484 46954 2484 46954 0 net4
rlabel metal1 2116 57426 2116 57426 0 net40
rlabel metal1 58282 24786 58282 24786 0 net41
rlabel metal2 53130 4454 53130 4454 0 net42
rlabel metal1 32246 13498 32246 13498 0 net43
rlabel metal1 39192 7990 39192 7990 0 net44
rlabel metal1 36064 18054 36064 18054 0 net45
rlabel metal1 35006 2550 35006 2550 0 net46
rlabel metal1 46651 3094 46651 3094 0 net47
rlabel metal1 40296 2482 40296 2482 0 net48
rlabel metal1 35006 4488 35006 4488 0 net49
rlabel metal1 57178 25194 57178 25194 0 net5
rlabel metal1 58144 22202 58144 22202 0 net6
rlabel metal1 57638 24378 57638 24378 0 net7
rlabel metal1 4508 57426 4508 57426 0 net8
rlabel metal1 2162 53550 2162 53550 0 net9
rlabel metal2 44482 20383 44482 20383 0 p_shaping_I.bit_in
rlabel metal1 51934 19482 51934 19482 0 p_shaping_I.bit_in_1
rlabel metal1 45816 21998 45816 21998 0 p_shaping_I.bit_in_2
rlabel metal2 43470 23528 43470 23528 0 p_shaping_I.counter\[0\]
rlabel metal1 44068 23698 44068 23698 0 p_shaping_I.counter\[1\]
rlabel metal1 44068 19686 44068 19686 0 p_shaping_I.ctl_1
rlabel metal2 23782 16422 23782 16422 0 p_shaping_Q.bit_in_1
rlabel metal1 23920 16762 23920 16762 0 p_shaping_Q.bit_in_2
rlabel metal1 24104 19482 24104 19482 0 p_shaping_Q.counter\[0\]
rlabel metal1 27600 18258 27600 18258 0 p_shaping_Q.counter\[1\]
rlabel metal1 24564 14246 24564 14246 0 p_shaping_Q.ctl_1
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
