magic
tech sky130A
magscale 1 2
timestamp 1671750302
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 14 2128 58880 57712
<< metal2 >>
rect 6458 59200 6514 59800
rect 28354 59200 28410 59800
rect 49606 59200 49662 59800
rect 18 200 74 800
rect 21270 200 21326 800
rect 42522 200 42578 800
<< obsm2 >>
rect 20 59144 6402 59200
rect 6570 59144 28298 59200
rect 28466 59144 49550 59200
rect 49718 59144 58310 59200
rect 20 856 58310 59144
rect 130 800 21214 856
rect 21382 800 42466 856
rect 42634 800 58310 856
<< metal3 >>
rect 59200 48968 59800 49088
rect 200 44888 800 45008
rect 59200 26528 59800 26648
rect 200 22448 800 22568
rect 59200 3408 59800 3528
<< obsm3 >>
rect 800 49168 59200 57697
rect 800 48888 59120 49168
rect 800 45088 59200 48888
rect 880 44808 59200 45088
rect 800 26728 59200 44808
rect 800 26448 59120 26728
rect 800 22648 59200 26448
rect 880 22368 59200 22648
rect 800 3608 59200 22368
rect 800 3328 59120 3608
rect 800 2143 59200 3328
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< labels >>
rlabel metal3 s 200 44888 800 45008 6 clk
port 1 nsew signal input
rlabel metal3 s 59200 3408 59800 3528 6 cout1
port 2 nsew signal output
rlabel metal2 s 18 200 74 800 6 cout10
port 3 nsew signal output
rlabel metal2 s 49606 59200 49662 59800 6 cout2
port 4 nsew signal output
rlabel metal2 s 42522 200 42578 800 6 cout3
port 5 nsew signal output
rlabel metal3 s 200 22448 800 22568 6 cout4
port 6 nsew signal output
rlabel metal3 s 59200 48968 59800 49088 6 cout5
port 7 nsew signal output
rlabel metal2 s 21270 200 21326 800 6 cout6
port 8 nsew signal output
rlabel metal2 s 6458 59200 6514 59800 6 cout7
port 9 nsew signal output
rlabel metal2 s 28354 59200 28410 59800 6 cout8
port 10 nsew signal output
rlabel metal3 s 59200 26528 59800 26648 6 cout9
port 11 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2415526
string GDS_FILE /home/urielcho/Proyectos_caravel/MPW8/gf180_vs_sky130/openlane/divider/runs/22_12_22_17_03/results/signoff/divider.magic.gds
string GDS_START 247274
<< end >>

