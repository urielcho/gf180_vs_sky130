// This is the unpowered netlist.
module OQPSK_PS_RCOSINE2 (BitIn,
    CLK,
    EN,
    RST,
    I,
    Q,
    addI,
    addQ);
 input BitIn;
 input CLK;
 input EN;
 input RST;
 output [12:0] I;
 output [12:0] Q;
 output [5:0] addI;
 output [5:0] addQ;

 wire \Reg_Delay_Q.In ;
 wire \Reg_Delay_Q.Out ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire \bit2symb.regi ;
 wire \p_shaping_I.bit_in ;
 wire \p_shaping_I.bit_in_1 ;
 wire \p_shaping_I.bit_in_2 ;
 wire \p_shaping_I.counter[0] ;
 wire \p_shaping_I.counter[1] ;
 wire \p_shaping_I.ctl_1 ;
 wire \p_shaping_Q.bit_in_1 ;
 wire \p_shaping_Q.bit_in_2 ;
 wire \p_shaping_Q.counter[0] ;
 wire \p_shaping_Q.counter[1] ;
 wire \p_shaping_Q.ctl_1 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire clknet_0_CLK;
 wire clknet_1_0__leaf_CLK;
 wire clknet_1_1__leaf_CLK;

 sky130_fd_sc_hd__inv_2 _0985_ (.A(net33),
    .Y(_0803_));
 sky130_fd_sc_hd__and3_2 _0986_ (.A(net31),
    .B(net30),
    .C(net32),
    .X(_0814_));
 sky130_fd_sc_hd__clkbuf_4 _0987_ (.A(net32),
    .X(_0825_));
 sky130_fd_sc_hd__and2b_1 _0988_ (.A_N(_0825_),
    .B(net33),
    .X(_0835_));
 sky130_fd_sc_hd__a21oi_2 _0989_ (.A1(_0803_),
    .A2(_0814_),
    .B1(_0835_),
    .Y(_0846_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(net35),
    .Y(_0857_));
 sky130_fd_sc_hd__nor2_4 _0991_ (.A(_0857_),
    .B(net34),
    .Y(_0868_));
 sky130_fd_sc_hd__buf_2 _0992_ (.A(net31),
    .X(_0878_));
 sky130_fd_sc_hd__clkbuf_4 _0993_ (.A(net33),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_4 _0994_ (.A(net30),
    .X(_0900_));
 sky130_fd_sc_hd__or4b_4 _0995_ (.A(_0878_),
    .B(_0889_),
    .C(_0825_),
    .D_N(_0900_),
    .X(_0910_));
 sky130_fd_sc_hd__or2_1 _0996_ (.A(net31),
    .B(net32),
    .X(_0921_));
 sky130_fd_sc_hd__buf_2 _0997_ (.A(_0921_),
    .X(_0932_));
 sky130_fd_sc_hd__o211a_2 _0998_ (.A1(_0889_),
    .A2(_0932_),
    .B1(net34),
    .C1(net35),
    .X(_0942_));
 sky130_fd_sc_hd__a31oi_4 _0999_ (.A1(_0889_),
    .A2(net34),
    .A3(_0932_),
    .B1(net35),
    .Y(_0953_));
 sky130_fd_sc_hd__a2111oi_4 _1000_ (.A1(_0846_),
    .A2(_0868_),
    .B1(_0910_),
    .C1(_0942_),
    .D1(_0953_),
    .Y(_0004_));
 sky130_fd_sc_hd__clkbuf_4 _1001_ (.A(net37),
    .X(_0973_));
 sky130_fd_sc_hd__buf_2 _1002_ (.A(net39),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_4 _1003_ (.A(net44),
    .X(_0036_));
 sky130_fd_sc_hd__buf_4 _1004_ (.A(net36),
    .X(_0046_));
 sky130_fd_sc_hd__or4b_2 _1005_ (.A(_0973_),
    .B(_0984_),
    .C(_0036_),
    .D_N(_0046_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_4 _1006_ (.A(net44),
    .X(_0067_));
 sky130_fd_sc_hd__nand2_1 _1007_ (.A(_0984_),
    .B(_0067_),
    .Y(_0077_));
 sky130_fd_sc_hd__buf_2 _1008_ (.A(net37),
    .X(_0084_));
 sky130_fd_sc_hd__a31o_2 _1009_ (.A1(_0084_),
    .A2(_0046_),
    .A3(_0067_),
    .B1(_0984_),
    .X(_0090_));
 sky130_fd_sc_hd__or2b_1 _1010_ (.A(net43),
    .B_N(net41),
    .X(_0096_));
 sky130_fd_sc_hd__buf_2 _1011_ (.A(_0096_),
    .X(_0103_));
 sky130_fd_sc_hd__a21oi_1 _1012_ (.A1(_0077_),
    .A2(_0090_),
    .B1(_0103_),
    .Y(_0105_));
 sky130_fd_sc_hd__clkbuf_4 _1013_ (.A(_0984_),
    .X(_0106_));
 sky130_fd_sc_hd__or2_2 _1014_ (.A(_0973_),
    .B(net44),
    .X(_0107_));
 sky130_fd_sc_hd__o211a_1 _1015_ (.A1(_0106_),
    .A2(_0107_),
    .B1(net41),
    .C1(net43),
    .X(_0108_));
 sky130_fd_sc_hd__clkinv_2 _1016_ (.A(net43),
    .Y(_0109_));
 sky130_fd_sc_hd__o21ai_2 _1017_ (.A1(_0084_),
    .A2(_0067_),
    .B1(_0984_),
    .Y(_0110_));
 sky130_fd_sc_hd__clkinv_2 _1018_ (.A(net41),
    .Y(_0111_));
 sky130_fd_sc_hd__o21a_1 _1019_ (.A1(_0109_),
    .A2(_0110_),
    .B1(_0111_),
    .X(_0112_));
 sky130_fd_sc_hd__or4_4 _1020_ (.A(_0057_),
    .B(_0105_),
    .C(_0108_),
    .D(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__inv_2 _1021_ (.A(_0113_),
    .Y(_0005_));
 sky130_fd_sc_hd__clkbuf_4 _1022_ (.A(\p_shaping_I.bit_in ),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _1023_ (.A0(_0114_),
    .A1(\p_shaping_I.ctl_1 ),
    .S(net48),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(_0115_),
    .A1(\p_shaping_I.bit_in_1 ),
    .S(net42),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _1025_ (.A(_0116_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_2 _1026_ (.A(\p_shaping_Q.bit_in_1 ),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _1027_ (.A0(net45),
    .A1(\p_shaping_Q.ctl_1 ),
    .S(net49),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _1028_ (.A0(_0117_),
    .A1(_0118_),
    .S(_0113_),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_1 _1029_ (.A(_0119_),
    .X(_0002_));
 sky130_fd_sc_hd__and2b_1 _1030_ (.A_N(_0004_),
    .B(net48),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _1031_ (.A(_0120_),
    .X(_0001_));
 sky130_fd_sc_hd__and2_1 _1032_ (.A(net49),
    .B(_0113_),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_1 _1033_ (.A(_0121_),
    .X(_0003_));
 sky130_fd_sc_hd__clkbuf_4 _1034_ (.A(_0111_),
    .X(_0122_));
 sky130_fd_sc_hd__buf_2 _1035_ (.A(_0109_),
    .X(_0123_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(net39),
    .Y(_0124_));
 sky130_fd_sc_hd__clkbuf_4 _1037_ (.A(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__buf_2 _1038_ (.A(net36),
    .X(_0126_));
 sky130_fd_sc_hd__nor2_2 _1039_ (.A(_0126_),
    .B(_0036_),
    .Y(_0127_));
 sky130_fd_sc_hd__or2_2 _1040_ (.A(_0125_),
    .B(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__buf_2 _1041_ (.A(_0973_),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_4 _1042_ (.A(_0126_),
    .X(_0130_));
 sky130_fd_sc_hd__nand2_1 _1043_ (.A(_0129_),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__or2b_1 _1044_ (.A(_0084_),
    .B_N(_0036_),
    .X(_0132_));
 sky130_fd_sc_hd__o21a_1 _1045_ (.A1(_0046_),
    .A2(_0067_),
    .B1(_0106_),
    .X(_0133_));
 sky130_fd_sc_hd__and3_1 _1046_ (.A(_0131_),
    .B(_0132_),
    .C(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_4 _1047_ (.A(_0036_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_4 _1048_ (.A(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__and2b_2 _1049_ (.A_N(_0126_),
    .B(net37),
    .X(_0137_));
 sky130_fd_sc_hd__nand2b_2 _1050_ (.A_N(_0126_),
    .B(net44),
    .Y(_0138_));
 sky130_fd_sc_hd__o211a_1 _1051_ (.A1(_0136_),
    .A2(_0137_),
    .B1(_0138_),
    .C1(_0125_),
    .X(_0139_));
 sky130_fd_sc_hd__a211o_1 _1052_ (.A1(_0123_),
    .A2(_0128_),
    .B1(_0134_),
    .C1(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__buf_2 _1053_ (.A(_0106_),
    .X(_0141_));
 sky130_fd_sc_hd__and2b_1 _1054_ (.A_N(_0973_),
    .B(net44),
    .X(_0142_));
 sky130_fd_sc_hd__nor2_1 _1055_ (.A(_0141_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(_0067_),
    .Y(_0144_));
 sky130_fd_sc_hd__xor2_4 _1057_ (.A(net37),
    .B(net36),
    .X(_0145_));
 sky130_fd_sc_hd__and3_1 _1058_ (.A(_0084_),
    .B(_0046_),
    .C(_0036_),
    .X(_0146_));
 sky130_fd_sc_hd__a211oi_2 _1059_ (.A1(_0144_),
    .A2(_0145_),
    .B1(_0146_),
    .C1(_0125_),
    .Y(_0147_));
 sky130_fd_sc_hd__and2b_1 _1060_ (.A_N(net43),
    .B(net41),
    .X(_0148_));
 sky130_fd_sc_hd__o21a_1 _1061_ (.A1(_0143_),
    .A2(_0147_),
    .B1(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__a211o_2 _1062_ (.A1(_0122_),
    .A2(_0140_),
    .B1(_0149_),
    .C1(_0108_),
    .X(_0150_));
 sky130_fd_sc_hd__nor2_4 _1063_ (.A(\p_shaping_Q.counter[1] ),
    .B(\p_shaping_Q.counter[0] ),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _1064_ (.A(\p_shaping_Q.counter[1] ),
    .Y(_0152_));
 sky130_fd_sc_hd__nor2_4 _1065_ (.A(_0973_),
    .B(_0046_),
    .Y(_0153_));
 sky130_fd_sc_hd__clkbuf_4 _1066_ (.A(_0106_),
    .X(_0154_));
 sky130_fd_sc_hd__a21oi_4 _1067_ (.A1(_0084_),
    .A2(_0046_),
    .B1(_0067_),
    .Y(_0155_));
 sky130_fd_sc_hd__nand2_2 _1068_ (.A(net43),
    .B(_0111_),
    .Y(_0156_));
 sky130_fd_sc_hd__nand2_1 _1069_ (.A(_0125_),
    .B(_0148_),
    .Y(_0157_));
 sky130_fd_sc_hd__o31a_1 _1070_ (.A1(_0154_),
    .A2(_0155_),
    .A3(_0156_),
    .B1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__or2_2 _1071_ (.A(net43),
    .B(net41),
    .X(_0159_));
 sky130_fd_sc_hd__a21oi_1 _1072_ (.A1(_0135_),
    .A2(_0145_),
    .B1(_0110_),
    .Y(_0160_));
 sky130_fd_sc_hd__o21a_1 _1073_ (.A1(_0135_),
    .A2(_0153_),
    .B1(_0124_),
    .X(_0161_));
 sky130_fd_sc_hd__a21bo_1 _1074_ (.A1(_0084_),
    .A2(_0067_),
    .B1_N(_0046_),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_1 _1075_ (.A(_0154_),
    .B(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__o32a_1 _1076_ (.A1(_0159_),
    .A2(_0160_),
    .A3(_0161_),
    .B1(_0156_),
    .B2(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__o21a_1 _1077_ (.A1(_0153_),
    .A2(_0158_),
    .B1(_0164_),
    .X(_0165_));
 sky130_fd_sc_hd__or2_2 _1078_ (.A(_0152_),
    .B(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(net37),
    .Y(_0167_));
 sky130_fd_sc_hd__and2b_1 _1080_ (.A_N(net44),
    .B(net36),
    .X(_0168_));
 sky130_fd_sc_hd__or4b_1 _1081_ (.A(_0167_),
    .B(_0106_),
    .C(_0168_),
    .D_N(_0138_),
    .X(_0169_));
 sky130_fd_sc_hd__a21bo_2 _1082_ (.A1(_0973_),
    .A2(_0036_),
    .B1_N(_0984_),
    .X(_0170_));
 sky130_fd_sc_hd__or2_1 _1083_ (.A(_0145_),
    .B(_0170_),
    .X(_0171_));
 sky130_fd_sc_hd__clkinv_2 _1084_ (.A(_0126_),
    .Y(_0172_));
 sky130_fd_sc_hd__a21o_2 _1085_ (.A1(_0084_),
    .A2(_0036_),
    .B1(_0984_),
    .X(_0173_));
 sky130_fd_sc_hd__o221a_1 _1086_ (.A1(_0172_),
    .A2(_0077_),
    .B1(_0153_),
    .B2(_0173_),
    .C1(net43),
    .X(_0174_));
 sky130_fd_sc_hd__a31o_1 _1087_ (.A1(_0109_),
    .A2(_0169_),
    .A3(_0171_),
    .B1(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__clkbuf_4 _1088_ (.A(net43),
    .X(_0176_));
 sky130_fd_sc_hd__nor2b_4 _1089_ (.A(_0036_),
    .B_N(_0973_),
    .Y(_0177_));
 sky130_fd_sc_hd__a21oi_1 _1090_ (.A1(_0125_),
    .A2(_0132_),
    .B1(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__or2b_1 _1091_ (.A(_0067_),
    .B_N(_0084_),
    .X(_0179_));
 sky130_fd_sc_hd__nor2_1 _1092_ (.A(_0106_),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__or4_4 _1093_ (.A(net37),
    .B(_0126_),
    .C(net39),
    .D(net44),
    .X(_0181_));
 sky130_fd_sc_hd__o311a_1 _1094_ (.A1(_0176_),
    .A2(_0178_),
    .A3(_0180_),
    .B1(_0181_),
    .C1(net41),
    .X(_0182_));
 sky130_fd_sc_hd__a21o_2 _1095_ (.A1(_0122_),
    .A2(_0175_),
    .B1(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__xnor2_2 _1096_ (.A(_0166_),
    .B(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__nor2_1 _1097_ (.A(_0151_),
    .B(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__xnor2_2 _1098_ (.A(_0150_),
    .B(_0185_),
    .Y(net17));
 sky130_fd_sc_hd__inv_2 _1099_ (.A(_0151_),
    .Y(_0186_));
 sky130_fd_sc_hd__buf_2 _1100_ (.A(_0186_),
    .X(_0022_));
 sky130_fd_sc_hd__buf_2 _1101_ (.A(\p_shaping_Q.bit_in_2 ),
    .X(_0187_));
 sky130_fd_sc_hd__clkbuf_4 _1102_ (.A(net41),
    .X(_0188_));
 sky130_fd_sc_hd__a21oi_4 _1103_ (.A1(_0067_),
    .A2(_0145_),
    .B1(_0106_),
    .Y(_0189_));
 sky130_fd_sc_hd__a211o_1 _1104_ (.A1(_0132_),
    .A2(_0133_),
    .B1(_0189_),
    .C1(_0176_),
    .X(_0190_));
 sky130_fd_sc_hd__xnor2_4 _1105_ (.A(_0973_),
    .B(_0046_),
    .Y(_0191_));
 sky130_fd_sc_hd__nor2_1 _1106_ (.A(_0125_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__and2b_1 _1107_ (.A_N(_0973_),
    .B(_0126_),
    .X(_0193_));
 sky130_fd_sc_hd__or4bb_1 _1108_ (.A(net37),
    .B(_0126_),
    .C_N(_0984_),
    .D_N(net44),
    .X(_0194_));
 sky130_fd_sc_hd__o31a_1 _1109_ (.A1(_0106_),
    .A2(_0135_),
    .A3(_0193_),
    .B1(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__a21o_1 _1110_ (.A1(net43),
    .A2(_0181_),
    .B1(_0111_),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _1111_ (.A(_0195_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__o221a_1 _1112_ (.A1(_0188_),
    .A2(_0190_),
    .B1(_0192_),
    .B2(_0156_),
    .C1(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__and2_1 _1113_ (.A(_0165_),
    .B(_0198_),
    .X(_0199_));
 sky130_fd_sc_hd__and2b_1 _1114_ (.A_N(_0984_),
    .B(_0036_),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_2 _1115_ (.A(_0130_),
    .B(_0067_),
    .Y(_0201_));
 sky130_fd_sc_hd__o21a_1 _1116_ (.A1(_0154_),
    .A2(_0137_),
    .B1(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__nand2_2 _1117_ (.A(_0125_),
    .B(_0201_),
    .Y(_0203_));
 sky130_fd_sc_hd__and3b_2 _1118_ (.A_N(net37),
    .B(_0126_),
    .C(net44),
    .X(_0204_));
 sky130_fd_sc_hd__a2111oi_1 _1119_ (.A1(_0154_),
    .A2(_0204_),
    .B1(_0127_),
    .C1(_0177_),
    .D1(_0176_),
    .Y(_0205_));
 sky130_fd_sc_hd__and3b_1 _1120_ (.A_N(_0036_),
    .B(_0046_),
    .C(_0084_),
    .X(_0206_));
 sky130_fd_sc_hd__a21o_1 _1121_ (.A1(_0125_),
    .A2(_0206_),
    .B1(_0109_),
    .X(_0207_));
 sky130_fd_sc_hd__o32a_1 _1122_ (.A1(_0106_),
    .A2(_0135_),
    .A3(_0193_),
    .B1(_0155_),
    .B2(_0146_),
    .X(_0208_));
 sky130_fd_sc_hd__o2bb2a_1 _1123_ (.A1_N(_0203_),
    .A2_N(_0205_),
    .B1(_0207_),
    .B2(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__o32a_1 _1124_ (.A1(_0103_),
    .A2(_0200_),
    .A3(_0202_),
    .B1(_0209_),
    .B2(_0188_),
    .X(_0210_));
 sky130_fd_sc_hd__or3_1 _1125_ (.A(_0187_),
    .B(_0199_),
    .C(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__o21ai_1 _1126_ (.A1(_0187_),
    .A2(_0199_),
    .B1(_0210_),
    .Y(_0212_));
 sky130_fd_sc_hd__or2b_2 _1127_ (.A(_0046_),
    .B_N(_0084_),
    .X(_0213_));
 sky130_fd_sc_hd__o211ai_4 _1128_ (.A1(_0135_),
    .A2(_0213_),
    .B1(_0201_),
    .C1(_0154_),
    .Y(_0214_));
 sky130_fd_sc_hd__o31a_1 _1129_ (.A1(_0130_),
    .A2(_0142_),
    .A3(_0177_),
    .B1(_0109_),
    .X(_0215_));
 sky130_fd_sc_hd__and4_1 _1130_ (.A(_0973_),
    .B(_0126_),
    .C(_0984_),
    .D(net44),
    .X(_0216_));
 sky130_fd_sc_hd__and2_1 _1131_ (.A(net43),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__a211o_1 _1132_ (.A1(_0214_),
    .A2(_0215_),
    .B1(_0217_),
    .C1(_0180_),
    .X(_0218_));
 sky130_fd_sc_hd__nor2_1 _1133_ (.A(_0135_),
    .B(_0145_),
    .Y(_0219_));
 sky130_fd_sc_hd__o221a_1 _1134_ (.A1(_0135_),
    .A2(_0191_),
    .B1(_0138_),
    .B2(_0129_),
    .C1(_0154_),
    .X(_0220_));
 sky130_fd_sc_hd__nor4_1 _1135_ (.A(_0176_),
    .B(_0204_),
    .C(_0219_),
    .D(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__o31a_1 _1136_ (.A1(_0154_),
    .A2(_0111_),
    .A3(_0107_),
    .B1(_0103_),
    .X(_0222_));
 sky130_fd_sc_hd__o2bb2a_1 _1137_ (.A1_N(_0122_),
    .A2_N(_0218_),
    .B1(_0221_),
    .B2(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__a211o_1 _1138_ (.A1(_0122_),
    .A2(_0175_),
    .B1(_0182_),
    .C1(\p_shaping_Q.bit_in_1 ),
    .X(_0224_));
 sky130_fd_sc_hd__o21a_1 _1139_ (.A1(_0117_),
    .A2(_0223_),
    .B1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__o21bai_2 _1140_ (.A1(_0130_),
    .A2(_0135_),
    .B1_N(_0129_),
    .Y(_0226_));
 sky130_fd_sc_hd__and2_1 _1141_ (.A(_0154_),
    .B(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__a21o_1 _1142_ (.A1(_0176_),
    .A2(_0057_),
    .B1(_0111_),
    .X(_0228_));
 sky130_fd_sc_hd__o21bai_1 _1143_ (.A1(_0189_),
    .A2(_0227_),
    .B1_N(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__a2bb2o_1 _1144_ (.A1_N(_0130_),
    .A2_N(_0170_),
    .B1(_0137_),
    .B2(_0200_),
    .X(_0230_));
 sky130_fd_sc_hd__or4_2 _1145_ (.A(_0106_),
    .B(_0137_),
    .C(_0127_),
    .D(_0204_),
    .X(_0231_));
 sky130_fd_sc_hd__a21oi_1 _1146_ (.A1(_0154_),
    .A2(_0226_),
    .B1(_0176_),
    .Y(_0232_));
 sky130_fd_sc_hd__a221o_1 _1147_ (.A1(_0176_),
    .A2(_0230_),
    .B1(_0231_),
    .B2(_0232_),
    .C1(net41),
    .X(_0233_));
 sky130_fd_sc_hd__and2_1 _1148_ (.A(_0229_),
    .B(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__a21oi_1 _1149_ (.A1(net49),
    .A2(\p_shaping_Q.ctl_1 ),
    .B1(net45),
    .Y(_0235_));
 sky130_fd_sc_hd__and3_1 _1150_ (.A(net49),
    .B(net45),
    .C(\p_shaping_Q.ctl_1 ),
    .X(_0236_));
 sky130_fd_sc_hd__nor3_2 _1151_ (.A(_0113_),
    .B(_0235_),
    .C(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__nor2_1 _1152_ (.A(_0234_),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__xnor2_1 _1153_ (.A(_0225_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__a31o_1 _1154_ (.A1(\p_shaping_Q.counter[1] ),
    .A2(_0211_),
    .A3(_0212_),
    .B1(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__buf_2 _1155_ (.A(\p_shaping_Q.counter[1] ),
    .X(_0241_));
 sky130_fd_sc_hd__nand4_1 _1156_ (.A(_0241_),
    .B(_0211_),
    .C(_0212_),
    .D(_0239_),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _1157_ (.A(net45),
    .Y(_0243_));
 sky130_fd_sc_hd__buf_2 _1158_ (.A(_0125_),
    .X(_0244_));
 sky130_fd_sc_hd__mux4_1 _1159_ (.A0(_0107_),
    .A1(_0146_),
    .A2(_0226_),
    .A3(_0137_),
    .S0(_0109_),
    .S1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__buf_2 _1160_ (.A(_0176_),
    .X(_0246_));
 sky130_fd_sc_hd__nor2_1 _1161_ (.A(_0167_),
    .B(_0172_),
    .Y(_0247_));
 sky130_fd_sc_hd__o41a_1 _1162_ (.A1(_0136_),
    .A2(_0246_),
    .A3(_0247_),
    .A4(_0133_),
    .B1(_0188_),
    .X(_0248_));
 sky130_fd_sc_hd__a2bb2o_2 _1163_ (.A1_N(_0188_),
    .A2_N(_0245_),
    .B1(_0190_),
    .B2(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_1 _1164_ (.A(_0150_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__and2_1 _1165_ (.A(_0243_),
    .B(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__a21oi_2 _1166_ (.A1(_0141_),
    .A2(_0144_),
    .B1(_0246_),
    .Y(_0252_));
 sky130_fd_sc_hd__nand2_1 _1167_ (.A(_0141_),
    .B(_0131_),
    .Y(_0253_));
 sky130_fd_sc_hd__or3_1 _1168_ (.A(_0154_),
    .B(_0204_),
    .C(_0206_),
    .X(_0254_));
 sky130_fd_sc_hd__a21boi_1 _1169_ (.A1(_0129_),
    .A2(_0130_),
    .B1_N(_0135_),
    .Y(_0255_));
 sky130_fd_sc_hd__o221a_1 _1170_ (.A1(_0136_),
    .A2(_0145_),
    .B1(_0255_),
    .B2(_0125_),
    .C1(_0176_),
    .X(_0256_));
 sky130_fd_sc_hd__a31o_1 _1171_ (.A1(_0252_),
    .A2(_0253_),
    .A3(_0254_),
    .B1(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__buf_2 _1172_ (.A(_0141_),
    .X(_0258_));
 sky130_fd_sc_hd__o311a_1 _1173_ (.A1(_0172_),
    .A2(_0258_),
    .A3(_0177_),
    .B1(_0163_),
    .C1(_0148_),
    .X(_0259_));
 sky130_fd_sc_hd__a21oi_2 _1174_ (.A1(_0122_),
    .A2(_0257_),
    .B1(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__xnor2_1 _1175_ (.A(_0251_),
    .B(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand4_1 _1176_ (.A(_0022_),
    .B(_0240_),
    .C(_0242_),
    .D(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__a31o_1 _1177_ (.A1(_0186_),
    .A2(_0240_),
    .A3(_0242_),
    .B1(_0261_),
    .X(_0263_));
 sky130_fd_sc_hd__o21ai_1 _1178_ (.A1(\p_shaping_Q.bit_in_2 ),
    .A2(_0165_),
    .B1(_0198_),
    .Y(_0264_));
 sky130_fd_sc_hd__or3_1 _1179_ (.A(\p_shaping_Q.bit_in_2 ),
    .B(_0165_),
    .C(_0198_),
    .X(_0265_));
 sky130_fd_sc_hd__xor2_1 _1180_ (.A(_0224_),
    .B(_0223_),
    .X(_0266_));
 sky130_fd_sc_hd__a31o_1 _1181_ (.A1(\p_shaping_Q.counter[1] ),
    .A2(_0264_),
    .A3(_0265_),
    .B1(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__nor2_1 _1182_ (.A(net45),
    .B(_0150_),
    .Y(_0268_));
 sky130_fd_sc_hd__xnor2_2 _1183_ (.A(_0249_),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__and4_1 _1184_ (.A(\p_shaping_Q.counter[1] ),
    .B(_0264_),
    .C(_0265_),
    .D(_0266_),
    .X(_0270_));
 sky130_fd_sc_hd__a31o_1 _1185_ (.A1(_0186_),
    .A2(_0267_),
    .A3(_0269_),
    .B1(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__a21oi_1 _1186_ (.A1(_0262_),
    .A2(_0263_),
    .B1(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__and3_1 _1187_ (.A(_0262_),
    .B(_0263_),
    .C(_0271_),
    .X(_0273_));
 sky130_fd_sc_hd__or2_1 _1188_ (.A(_0272_),
    .B(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__or3b_1 _1189_ (.A(_0151_),
    .B(_0270_),
    .C_N(_0267_),
    .X(_0275_));
 sky130_fd_sc_hd__xor2_2 _1190_ (.A(_0275_),
    .B(_0269_),
    .X(_0276_));
 sky130_fd_sc_hd__o32ai_4 _1191_ (.A1(_0150_),
    .A2(_0151_),
    .A3(_0184_),
    .B1(_0166_),
    .B2(_0183_),
    .Y(_0277_));
 sky130_fd_sc_hd__and2b_1 _1192_ (.A_N(_0276_),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__xnor2_2 _1193_ (.A(_0274_),
    .B(_0278_),
    .Y(net22));
 sky130_fd_sc_hd__and4_1 _1194_ (.A(_0241_),
    .B(_0211_),
    .C(_0212_),
    .D(_0239_),
    .X(_0279_));
 sky130_fd_sc_hd__and4_1 _1195_ (.A(_0022_),
    .B(_0240_),
    .C(_0242_),
    .D(_0261_),
    .X(_0280_));
 sky130_fd_sc_hd__and3_1 _1196_ (.A(_0165_),
    .B(_0198_),
    .C(_0210_),
    .X(_0281_));
 sky130_fd_sc_hd__nor2_1 _1197_ (.A(_0141_),
    .B(_0153_),
    .Y(_0282_));
 sky130_fd_sc_hd__a21o_1 _1198_ (.A1(_0136_),
    .A2(_0213_),
    .B1(_0177_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _1199_ (.A0(_0258_),
    .A1(_0282_),
    .S(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__nor2_1 _1200_ (.A(_0146_),
    .B(_0155_),
    .Y(_0285_));
 sky130_fd_sc_hd__or2_1 _1201_ (.A(_0168_),
    .B(_0173_),
    .X(_0286_));
 sky130_fd_sc_hd__nor2_1 _1202_ (.A(_0246_),
    .B(_0188_),
    .Y(_0287_));
 sky130_fd_sc_hd__o211ai_1 _1203_ (.A1(_0128_),
    .A2(_0285_),
    .B1(_0286_),
    .C1(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _1204_ (.A(_0244_),
    .B(_0226_),
    .Y(_0289_));
 sky130_fd_sc_hd__a21o_1 _1205_ (.A1(_0136_),
    .A2(_0191_),
    .B1(_0127_),
    .X(_0290_));
 sky130_fd_sc_hd__a21oi_1 _1206_ (.A1(_0289_),
    .A2(_0290_),
    .B1(_0103_),
    .Y(_0291_));
 sky130_fd_sc_hd__o21ai_1 _1207_ (.A1(_0289_),
    .A2(_0290_),
    .B1(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__o211a_1 _1208_ (.A1(_0156_),
    .A2(_0284_),
    .B1(_0288_),
    .C1(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__o21ai_1 _1209_ (.A1(_0187_),
    .A2(_0281_),
    .B1(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__or3_1 _1210_ (.A(_0187_),
    .B(_0293_),
    .C(_0281_),
    .X(_0295_));
 sky130_fd_sc_hd__a31o_1 _1211_ (.A1(_0183_),
    .A2(_0223_),
    .A3(_0234_),
    .B1(_0117_),
    .X(_0296_));
 sky130_fd_sc_hd__nor2_1 _1212_ (.A(_0143_),
    .B(_0220_),
    .Y(_0297_));
 sky130_fd_sc_hd__a211oi_1 _1213_ (.A1(_0244_),
    .A2(_0283_),
    .B1(_0160_),
    .C1(_0246_),
    .Y(_0298_));
 sky130_fd_sc_hd__a31o_1 _1214_ (.A1(_0246_),
    .A2(_0203_),
    .A3(_0163_),
    .B1(_0188_),
    .X(_0299_));
 sky130_fd_sc_hd__o22ai_2 _1215_ (.A1(_0196_),
    .A2(_0297_),
    .B1(_0298_),
    .B2(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__or2_1 _1216_ (.A(_0237_),
    .B(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__xnor2_1 _1217_ (.A(_0296_),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__a31o_1 _1218_ (.A1(\p_shaping_Q.counter[1] ),
    .A2(_0294_),
    .A3(_0295_),
    .B1(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__nand4_1 _1219_ (.A(_0241_),
    .B(_0294_),
    .C(_0295_),
    .D(_0302_),
    .Y(_0304_));
 sky130_fd_sc_hd__and3_1 _1220_ (.A(_0186_),
    .B(_0303_),
    .C(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__a31o_1 _1221_ (.A1(_0150_),
    .A2(_0249_),
    .A3(_0260_),
    .B1(net45),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_1 _1222_ (.A(_0144_),
    .B(_0191_),
    .Y(_0307_));
 sky130_fd_sc_hd__o221a_1 _1223_ (.A1(_0191_),
    .A2(_0128_),
    .B1(_0307_),
    .B2(_0258_),
    .C1(_0148_),
    .X(_0308_));
 sky130_fd_sc_hd__o32a_1 _1224_ (.A1(_0130_),
    .A2(_0200_),
    .A3(_0177_),
    .B1(_0153_),
    .B2(_0258_),
    .X(_0309_));
 sky130_fd_sc_hd__nand2_1 _1225_ (.A(_0136_),
    .B(_0213_),
    .Y(_0310_));
 sky130_fd_sc_hd__and2_1 _1226_ (.A(_0141_),
    .B(_0162_),
    .X(_0311_));
 sky130_fd_sc_hd__a211o_1 _1227_ (.A1(_0244_),
    .A2(_0310_),
    .B1(_0311_),
    .C1(_0159_),
    .X(_0312_));
 sky130_fd_sc_hd__o221ai_1 _1228_ (.A1(_0122_),
    .A2(_0057_),
    .B1(_0156_),
    .B2(_0309_),
    .C1(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__or2_1 _1229_ (.A(_0308_),
    .B(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__xor2_1 _1230_ (.A(_0306_),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__xnor2_1 _1231_ (.A(_0305_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__o21a_1 _1232_ (.A1(_0279_),
    .A2(_0280_),
    .B1(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__or3_2 _1233_ (.A(_0279_),
    .B(_0280_),
    .C(_0316_),
    .X(_0318_));
 sky130_fd_sc_hd__and2b_1 _1234_ (.A_N(_0317_),
    .B(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _1235_ (.A1(_0262_),
    .A2(_0263_),
    .B1(_0271_),
    .X(_0320_));
 sky130_fd_sc_hd__a21o_2 _1236_ (.A1(_0320_),
    .A2(_0278_),
    .B1(_0273_),
    .X(_0321_));
 sky130_fd_sc_hd__xor2_2 _1237_ (.A(_0319_),
    .B(_0321_),
    .X(net23));
 sky130_fd_sc_hd__a21o_1 _1238_ (.A1(_0293_),
    .A2(_0281_),
    .B1(_0187_),
    .X(_0322_));
 sky130_fd_sc_hd__nor2_1 _1239_ (.A(_0145_),
    .B(_0170_),
    .Y(_0323_));
 sky130_fd_sc_hd__nor2_1 _1240_ (.A(_0323_),
    .B(_0189_),
    .Y(_0324_));
 sky130_fd_sc_hd__and2_1 _1241_ (.A(_0123_),
    .B(_0173_),
    .X(_0325_));
 sky130_fd_sc_hd__nor2_1 _1242_ (.A(_0167_),
    .B(_0168_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_2 _1243_ (.A(_0141_),
    .B(_0138_),
    .Y(_0327_));
 sky130_fd_sc_hd__o211a_1 _1244_ (.A1(_0326_),
    .A2(_0327_),
    .B1(_0231_),
    .C1(_0246_),
    .X(_0328_));
 sky130_fd_sc_hd__a21oi_1 _1245_ (.A1(_0253_),
    .A2(_0325_),
    .B1(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__o22a_1 _1246_ (.A1(_0103_),
    .A2(_0324_),
    .B1(_0329_),
    .B2(_0188_),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _1247_ (.A(_0322_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__or2_1 _1248_ (.A(_0322_),
    .B(_0330_),
    .X(_0332_));
 sky130_fd_sc_hd__inv_2 _1249_ (.A(_0117_),
    .Y(_0333_));
 sky130_fd_sc_hd__a21oi_1 _1250_ (.A1(_0229_),
    .A2(_0233_),
    .B1(_0117_),
    .Y(_0334_));
 sky130_fd_sc_hd__a21oi_1 _1251_ (.A1(_0333_),
    .A2(_0300_),
    .B1(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(_0225_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__o211a_1 _1253_ (.A1(_0129_),
    .A2(_0138_),
    .B1(_0179_),
    .C1(_0123_),
    .X(_0337_));
 sky130_fd_sc_hd__o31a_1 _1254_ (.A1(_0137_),
    .A2(_0128_),
    .A3(_0204_),
    .B1(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__nor2_1 _1255_ (.A(_0129_),
    .B(_0258_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _1256_ (.A(_0129_),
    .B(_0136_),
    .Y(_0340_));
 sky130_fd_sc_hd__and3_1 _1257_ (.A(_0258_),
    .B(_0107_),
    .C(_0340_),
    .X(_0341_));
 sky130_fd_sc_hd__a211o_1 _1258_ (.A1(_0172_),
    .A2(_0180_),
    .B1(_0193_),
    .C1(_0156_),
    .X(_0342_));
 sky130_fd_sc_hd__o31a_1 _1259_ (.A1(_0339_),
    .A2(_0159_),
    .A3(_0341_),
    .B1(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__or3_2 _1260_ (.A(_0113_),
    .B(_0235_),
    .C(_0236_),
    .X(_0344_));
 sky130_fd_sc_hd__o211a_1 _1261_ (.A1(_0196_),
    .A2(_0338_),
    .B1(_0343_),
    .C1(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__xnor2_1 _1262_ (.A(_0336_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__a31oi_1 _1263_ (.A1(_0241_),
    .A2(_0331_),
    .A3(_0332_),
    .B1(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__and4_1 _1264_ (.A(_0241_),
    .B(_0331_),
    .C(_0332_),
    .D(_0346_),
    .X(_0348_));
 sky130_fd_sc_hd__o31a_1 _1265_ (.A1(_0129_),
    .A2(_0244_),
    .A3(_0168_),
    .B1(_0203_),
    .X(_0349_));
 sky130_fd_sc_hd__a2bb2o_1 _1266_ (.A1_N(_0123_),
    .A2_N(_0349_),
    .B1(_0325_),
    .B2(_0129_),
    .X(_0350_));
 sky130_fd_sc_hd__nor2_1 _1267_ (.A(_0144_),
    .B(_0153_),
    .Y(_0351_));
 sky130_fd_sc_hd__nor2_1 _1268_ (.A(_0155_),
    .B(_0351_),
    .Y(_0352_));
 sky130_fd_sc_hd__or3_1 _1269_ (.A(_0141_),
    .B(_0247_),
    .C(_0127_),
    .X(_0353_));
 sky130_fd_sc_hd__o211a_1 _1270_ (.A1(_0244_),
    .A2(_0352_),
    .B1(_0353_),
    .C1(_0148_),
    .X(_0354_));
 sky130_fd_sc_hd__a21oi_1 _1271_ (.A1(_0122_),
    .A2(_0350_),
    .B1(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_2 _1272_ (.A(_0260_),
    .Y(_0356_));
 sky130_fd_sc_hd__o31a_1 _1273_ (.A1(_0250_),
    .A2(_0356_),
    .A3(_0314_),
    .B1(_0243_),
    .X(_0357_));
 sky130_fd_sc_hd__xor2_1 _1274_ (.A(_0355_),
    .B(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__or4_2 _1275_ (.A(_0151_),
    .B(_0347_),
    .C(_0348_),
    .D(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__o31ai_1 _1276_ (.A1(_0151_),
    .A2(_0347_),
    .A3(_0348_),
    .B1(_0358_),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _1277_ (.A(_0022_),
    .B(_0303_),
    .Y(_0361_));
 sky130_fd_sc_hd__o21ai_1 _1278_ (.A1(_0361_),
    .A2(_0315_),
    .B1(_0304_),
    .Y(_0362_));
 sky130_fd_sc_hd__a21o_1 _1279_ (.A1(_0359_),
    .A2(_0360_),
    .B1(_0362_),
    .X(_0363_));
 sky130_fd_sc_hd__nand3_2 _1280_ (.A(_0359_),
    .B(_0360_),
    .C(_0362_),
    .Y(_0364_));
 sky130_fd_sc_hd__o2111ai_4 _1281_ (.A1(_0317_),
    .A2(_0321_),
    .B1(_0363_),
    .C1(_0364_),
    .D1(_0318_),
    .Y(_0365_));
 sky130_fd_sc_hd__o21a_1 _1282_ (.A1(_0317_),
    .A2(_0321_),
    .B1(_0318_),
    .X(_0366_));
 sky130_fd_sc_hd__a21o_1 _1283_ (.A1(_0363_),
    .A2(_0364_),
    .B1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _1284_ (.A(_0365_),
    .B(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__clkbuf_1 _1285_ (.A(_0368_),
    .X(net24));
 sky130_fd_sc_hd__inv_2 _1286_ (.A(_0359_),
    .Y(_0369_));
 sky130_fd_sc_hd__or2_1 _1287_ (.A(_0244_),
    .B(_0155_),
    .X(_0370_));
 sky130_fd_sc_hd__nand2_1 _1288_ (.A(_0090_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__a21o_1 _1289_ (.A1(_0169_),
    .A2(_0327_),
    .B1(_0159_),
    .X(_0372_));
 sky130_fd_sc_hd__nor2_2 _1290_ (.A(_0123_),
    .B(_0188_),
    .Y(_0373_));
 sky130_fd_sc_hd__a31o_1 _1291_ (.A1(_0107_),
    .A2(_0340_),
    .A3(_0282_),
    .B1(_0323_),
    .X(_0374_));
 sky130_fd_sc_hd__nand2_1 _1292_ (.A(_0373_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__o211a_1 _1293_ (.A1(_0103_),
    .A2(_0371_),
    .B1(_0372_),
    .C1(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__a31o_1 _1294_ (.A1(_0293_),
    .A2(_0281_),
    .A3(_0330_),
    .B1(_0187_),
    .X(_0377_));
 sky130_fd_sc_hd__xor2_1 _1295_ (.A(_0376_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__or3_1 _1296_ (.A(_0141_),
    .B(_0137_),
    .C(_0204_),
    .X(_0379_));
 sky130_fd_sc_hd__o2bb2a_1 _1297_ (.A1_N(_0244_),
    .A2_N(_0155_),
    .B1(_0170_),
    .B2(_0130_),
    .X(_0380_));
 sky130_fd_sc_hd__a211o_1 _1298_ (.A1(_0379_),
    .A2(_0327_),
    .B1(_0380_),
    .C1(_0156_),
    .X(_0381_));
 sky130_fd_sc_hd__or4_1 _1299_ (.A(_0130_),
    .B(_0141_),
    .C(_0142_),
    .D(_0177_),
    .X(_0382_));
 sky130_fd_sc_hd__a21oi_1 _1300_ (.A1(_0258_),
    .A2(_0127_),
    .B1(_0103_),
    .Y(_0383_));
 sky130_fd_sc_hd__a22oi_1 _1301_ (.A1(_0287_),
    .A2(_0380_),
    .B1(_0382_),
    .B2(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__a21oi_1 _1302_ (.A1(_0381_),
    .A2(_0384_),
    .B1(_0117_),
    .Y(_0385_));
 sky130_fd_sc_hd__a31o_1 _1303_ (.A1(_0335_),
    .A2(_0381_),
    .A3(_0384_),
    .B1(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__a211o_2 _1304_ (.A1(_0333_),
    .A2(_0300_),
    .B1(_0385_),
    .C1(_0334_),
    .X(_0387_));
 sky130_fd_sc_hd__or2_1 _1305_ (.A(_0344_),
    .B(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__o21ai_1 _1306_ (.A1(_0237_),
    .A2(_0386_),
    .B1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__a21o_1 _1307_ (.A1(_0241_),
    .A2(_0378_),
    .B1(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__nand3_1 _1308_ (.A(_0241_),
    .B(_0378_),
    .C(_0389_),
    .Y(_0391_));
 sky130_fd_sc_hd__and3_1 _1309_ (.A(_0022_),
    .B(_0390_),
    .C(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__nor4b_1 _1310_ (.A(_0250_),
    .B(_0356_),
    .C(_0314_),
    .D_N(_0355_),
    .Y(_0393_));
 sky130_fd_sc_hd__or2_1 _1311_ (.A(\Reg_Delay_Q.Out ),
    .B(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__and2_1 _1312_ (.A(_0123_),
    .B(_0077_),
    .X(_0395_));
 sky130_fd_sc_hd__o21ai_1 _1313_ (.A1(_0203_),
    .A2(_0219_),
    .B1(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__a21oi_1 _1314_ (.A1(_0181_),
    .A2(_0396_),
    .B1(_0122_),
    .Y(_0397_));
 sky130_fd_sc_hd__buf_2 _1315_ (.A(_0258_),
    .X(_0398_));
 sky130_fd_sc_hd__and3_1 _1316_ (.A(_0398_),
    .B(_0144_),
    .C(_0287_),
    .X(_0399_));
 sky130_fd_sc_hd__a311oi_4 _1317_ (.A1(_0373_),
    .A2(_0173_),
    .A3(_0214_),
    .B1(_0397_),
    .C1(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__xnor2_1 _1318_ (.A(_0394_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__xnor2_1 _1319_ (.A(_0392_),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__o21a_1 _1320_ (.A1(_0348_),
    .A2(_0369_),
    .B1(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__nor3_1 _1321_ (.A(_0348_),
    .B(_0369_),
    .C(_0402_),
    .Y(_0404_));
 sky130_fd_sc_hd__nor2_2 _1322_ (.A(_0403_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__nand2_1 _1323_ (.A(_0364_),
    .B(_0365_),
    .Y(_0406_));
 sky130_fd_sc_hd__xor2_4 _1324_ (.A(_0405_),
    .B(_0406_),
    .X(net25));
 sky130_fd_sc_hd__inv_2 _1325_ (.A(_0187_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand4_2 _1326_ (.A(_0293_),
    .B(_0281_),
    .C(_0330_),
    .D(_0376_),
    .Y(_0408_));
 sky130_fd_sc_hd__nor2_1 _1327_ (.A(_0203_),
    .B(_0206_),
    .Y(_0409_));
 sky130_fd_sc_hd__and3_1 _1328_ (.A(_0258_),
    .B(_0123_),
    .C(_0142_),
    .X(_0410_));
 sky130_fd_sc_hd__nor2_1 _1329_ (.A(_0409_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__or2_1 _1330_ (.A(_0144_),
    .B(_0153_),
    .X(_0412_));
 sky130_fd_sc_hd__nand2_1 _1331_ (.A(_0144_),
    .B(_0153_),
    .Y(_0413_));
 sky130_fd_sc_hd__and3_1 _1332_ (.A(_0246_),
    .B(_0412_),
    .C(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _1333_ (.A0(_0411_),
    .A1(_0409_),
    .S(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__buf_2 _1334_ (.A(_0246_),
    .X(_0416_));
 sky130_fd_sc_hd__nor2_1 _1335_ (.A(_0416_),
    .B(_0090_),
    .Y(_0417_));
 sky130_fd_sc_hd__mux2_1 _1336_ (.A0(_0415_),
    .A1(_0417_),
    .S(_0188_),
    .X(_0418_));
 sky130_fd_sc_hd__a21o_1 _1337_ (.A1(_0407_),
    .A2(_0408_),
    .B1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__a31oi_1 _1338_ (.A1(_0407_),
    .A2(_0418_),
    .A3(_0408_),
    .B1(_0152_),
    .Y(_0420_));
 sky130_fd_sc_hd__buf_2 _1339_ (.A(_0188_),
    .X(_0421_));
 sky130_fd_sc_hd__o211a_1 _1340_ (.A1(_0136_),
    .A2(_0193_),
    .B1(_0412_),
    .C1(_0176_),
    .X(_0422_));
 sky130_fd_sc_hd__o21ai_1 _1341_ (.A1(_0398_),
    .A2(_0138_),
    .B1(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__or3_1 _1342_ (.A(_0258_),
    .B(_0138_),
    .C(_0422_),
    .X(_0424_));
 sky130_fd_sc_hd__o311a_1 _1343_ (.A1(_0246_),
    .A2(_0219_),
    .A3(_0327_),
    .B1(_0423_),
    .C1(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__xor2_1 _1344_ (.A(_0147_),
    .B(_0162_),
    .X(_0426_));
 sky130_fd_sc_hd__o221a_1 _1345_ (.A1(_0421_),
    .A2(_0425_),
    .B1(_0426_),
    .B2(_0103_),
    .C1(_0344_),
    .X(_0427_));
 sky130_fd_sc_hd__xnor2_1 _1346_ (.A(_0387_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__a21o_1 _1347_ (.A1(_0419_),
    .A2(_0420_),
    .B1(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__nand3_1 _1348_ (.A(_0419_),
    .B(_0420_),
    .C(_0428_),
    .Y(_0430_));
 sky130_fd_sc_hd__and3_2 _1349_ (.A(_0022_),
    .B(_0429_),
    .C(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__and2_1 _1350_ (.A(_0393_),
    .B(_0400_),
    .X(_0432_));
 sky130_fd_sc_hd__nor2_2 _1351_ (.A(net45),
    .B(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__a21o_1 _1352_ (.A1(_0136_),
    .A2(_0191_),
    .B1(_0110_),
    .X(_0434_));
 sky130_fd_sc_hd__a31o_1 _1353_ (.A1(_0416_),
    .A2(_0173_),
    .A3(_0434_),
    .B1(_0395_),
    .X(_0435_));
 sky130_fd_sc_hd__a21o_1 _1354_ (.A1(_0379_),
    .A2(_0327_),
    .B1(_0103_),
    .X(_0436_));
 sky130_fd_sc_hd__o21a_1 _1355_ (.A1(_0421_),
    .A2(_0435_),
    .B1(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__xnor2_2 _1356_ (.A(_0433_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__xor2_4 _1357_ (.A(_0431_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_1 _1358_ (.A(_0022_),
    .B(_0390_),
    .Y(_0440_));
 sky130_fd_sc_hd__o21ai_2 _1359_ (.A1(_0440_),
    .A2(_0401_),
    .B1(_0391_),
    .Y(_0441_));
 sky130_fd_sc_hd__xnor2_4 _1360_ (.A(_0439_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__o21ai_1 _1361_ (.A1(_0348_),
    .A2(_0369_),
    .B1(_0402_),
    .Y(_0443_));
 sky130_fd_sc_hd__a31o_1 _1362_ (.A1(_0364_),
    .A2(_0365_),
    .A3(_0443_),
    .B1(_0404_),
    .X(_0444_));
 sky130_fd_sc_hd__xor2_4 _1363_ (.A(_0442_),
    .B(_0444_),
    .X(net26));
 sky130_fd_sc_hd__a31o_1 _1364_ (.A1(_0398_),
    .A2(_0416_),
    .A3(_0413_),
    .B1(_0421_),
    .X(_0445_));
 sky130_fd_sc_hd__o21a_1 _1365_ (.A1(_0142_),
    .A2(_0206_),
    .B1(_0416_),
    .X(_0446_));
 sky130_fd_sc_hd__a211oi_1 _1366_ (.A1(_0252_),
    .A2(_0231_),
    .B1(_0445_),
    .C1(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__and3_1 _1367_ (.A(_0407_),
    .B(_0408_),
    .C(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__a21oi_1 _1368_ (.A1(_0407_),
    .A2(_0408_),
    .B1(_0447_),
    .Y(_0449_));
 sky130_fd_sc_hd__nor2_1 _1369_ (.A(_0339_),
    .B(_0160_),
    .Y(_0450_));
 sky130_fd_sc_hd__a221o_1 _1370_ (.A1(_0398_),
    .A2(_0310_),
    .B1(_0307_),
    .B2(_0189_),
    .C1(_0123_),
    .X(_0451_));
 sky130_fd_sc_hd__nor2_1 _1371_ (.A(_0144_),
    .B(_0191_),
    .Y(_0452_));
 sky130_fd_sc_hd__or3b_1 _1372_ (.A(_0244_),
    .B(_0452_),
    .C_N(_0413_),
    .X(_0453_));
 sky130_fd_sc_hd__a31o_1 _1373_ (.A1(_0122_),
    .A2(_0286_),
    .A3(_0453_),
    .B1(_0373_),
    .X(_0454_));
 sky130_fd_sc_hd__a2bb2o_1 _1374_ (.A1_N(_0228_),
    .A2_N(_0450_),
    .B1(_0451_),
    .B2(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _1375_ (.A0(_0387_),
    .A1(_0117_),
    .S(_0455_),
    .X(_0456_));
 sky130_fd_sc_hd__and2_1 _1376_ (.A(_0237_),
    .B(_0336_),
    .X(_0457_));
 sky130_fd_sc_hd__a21oi_1 _1377_ (.A1(_0344_),
    .A2(_0456_),
    .B1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__o31ai_1 _1378_ (.A1(_0152_),
    .A2(_0448_),
    .A3(_0449_),
    .B1(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__or4_1 _1379_ (.A(_0152_),
    .B(_0458_),
    .C(_0448_),
    .D(_0449_),
    .X(_0460_));
 sky130_fd_sc_hd__and3_1 _1380_ (.A(_0022_),
    .B(_0459_),
    .C(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__and2b_1 _1381_ (.A_N(_0155_),
    .B(_0417_),
    .X(_0462_));
 sky130_fd_sc_hd__or4_1 _1382_ (.A(_0123_),
    .B(_0421_),
    .C(_0110_),
    .D(_0351_),
    .X(_0463_));
 sky130_fd_sc_hd__o31a_1 _1383_ (.A1(_0228_),
    .A2(_0410_),
    .A3(_0462_),
    .B1(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__xnor2_1 _1384_ (.A(_0433_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__xor2_1 _1385_ (.A(_0461_),
    .B(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__a21bo_1 _1386_ (.A1(_0431_),
    .A2(_0438_),
    .B1_N(_0430_),
    .X(_0467_));
 sky130_fd_sc_hd__nand2_1 _1387_ (.A(_0466_),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _1388_ (.A(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__nor2_1 _1389_ (.A(_0466_),
    .B(_0467_),
    .Y(_0470_));
 sky130_fd_sc_hd__nor2_1 _1390_ (.A(_0469_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__and2_1 _1391_ (.A(_0439_),
    .B(_0441_),
    .X(_0472_));
 sky130_fd_sc_hd__inv_2 _1392_ (.A(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__a311o_1 _1393_ (.A1(_0364_),
    .A2(_0365_),
    .A3(_0443_),
    .B1(_0404_),
    .C1(_0442_),
    .X(_0474_));
 sky130_fd_sc_hd__nand2_1 _1394_ (.A(_0473_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__xor2_2 _1395_ (.A(_0471_),
    .B(_0475_),
    .X(net27));
 sky130_fd_sc_hd__or3_1 _1396_ (.A(_0398_),
    .B(_0168_),
    .C(_0153_),
    .X(_0476_));
 sky130_fd_sc_hd__and2_1 _1397_ (.A(_0416_),
    .B(_0181_),
    .X(_0477_));
 sky130_fd_sc_hd__a21oi_1 _1398_ (.A1(_0189_),
    .A2(_0307_),
    .B1(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__or3b_1 _1399_ (.A(_0246_),
    .B(_0128_),
    .C_N(_0310_),
    .X(_0479_));
 sky130_fd_sc_hd__o41a_1 _1400_ (.A1(_0398_),
    .A2(_0159_),
    .A3(_0177_),
    .A4(_0452_),
    .B1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__o21ai_1 _1401_ (.A1(_0122_),
    .A2(_0478_),
    .B1(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__a31o_1 _1402_ (.A1(_0373_),
    .A2(_0170_),
    .A3(_0476_),
    .B1(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _1403_ (.A0(_0117_),
    .A1(_0387_),
    .S(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__or2_1 _1404_ (.A(_0151_),
    .B(_0457_),
    .X(_0484_));
 sky130_fd_sc_hd__o21ba_1 _1405_ (.A1(_0237_),
    .A2(_0483_),
    .B1_N(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__nand2_1 _1406_ (.A(_0407_),
    .B(_0408_),
    .Y(_0486_));
 sky130_fd_sc_hd__or2_1 _1407_ (.A(_0398_),
    .B(_0255_),
    .X(_0487_));
 sky130_fd_sc_hd__o21a_1 _1408_ (.A1(_0487_),
    .A2(_0219_),
    .B1(_0252_),
    .X(_0488_));
 sky130_fd_sc_hd__and3_1 _1409_ (.A(_0244_),
    .B(_0416_),
    .C(_0155_),
    .X(_0489_));
 sky130_fd_sc_hd__or3_1 _1410_ (.A(_0445_),
    .B(_0488_),
    .C(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__o311a_1 _1411_ (.A1(_0187_),
    .A2(_0477_),
    .A3(_0338_),
    .B1(_0486_),
    .C1(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__o21ai_1 _1412_ (.A1(_0187_),
    .A2(_0490_),
    .B1(_0241_),
    .Y(_0492_));
 sky130_fd_sc_hd__nor2_1 _1413_ (.A(_0491_),
    .B(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__xnor2_1 _1414_ (.A(_0485_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__or2_1 _1415_ (.A(_0108_),
    .B(_0112_),
    .X(_0495_));
 sky130_fd_sc_hd__nor2_1 _1416_ (.A(_0105_),
    .B(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__o221a_1 _1417_ (.A1(_0167_),
    .A2(_0327_),
    .B1(_0352_),
    .B2(_0398_),
    .C1(_0123_),
    .X(_0497_));
 sky130_fd_sc_hd__and2b_1 _1418_ (.A_N(_0497_),
    .B(_0432_),
    .X(_0498_));
 sky130_fd_sc_hd__nor2_1 _1419_ (.A(_0496_),
    .B(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__mux2_1 _1420_ (.A0(_0496_),
    .A1(_0499_),
    .S(_0243_),
    .X(_0500_));
 sky130_fd_sc_hd__xnor2_1 _1421_ (.A(_0494_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__a21bo_1 _1422_ (.A1(_0461_),
    .A2(_0465_),
    .B1_N(_0460_),
    .X(_0502_));
 sky130_fd_sc_hd__xnor2_2 _1423_ (.A(_0501_),
    .B(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__a31o_1 _1424_ (.A1(_0473_),
    .A2(_0474_),
    .A3(_0468_),
    .B1(_0470_),
    .X(_0504_));
 sky130_fd_sc_hd__xor2_2 _1425_ (.A(_0503_),
    .B(_0504_),
    .X(net28));
 sky130_fd_sc_hd__nand2_1 _1426_ (.A(_0485_),
    .B(_0493_),
    .Y(_0505_));
 sky130_fd_sc_hd__or2b_1 _1427_ (.A(_0494_),
    .B_N(_0500_),
    .X(_0506_));
 sky130_fd_sc_hd__a21o_1 _1428_ (.A1(_0144_),
    .A2(_0145_),
    .B1(_0170_),
    .X(_0507_));
 sky130_fd_sc_hd__a21o_1 _1429_ (.A1(_0487_),
    .A2(_0507_),
    .B1(_0416_),
    .X(_0508_));
 sky130_fd_sc_hd__nor2_1 _1430_ (.A(_0421_),
    .B(_0489_),
    .Y(_0509_));
 sky130_fd_sc_hd__a22o_1 _1431_ (.A1(_0421_),
    .A2(_0497_),
    .B1(_0508_),
    .B2(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(_0387_),
    .A1(_0117_),
    .S(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__o21bai_1 _1433_ (.A1(_0237_),
    .A2(_0511_),
    .B1_N(_0484_),
    .Y(_0512_));
 sky130_fd_sc_hd__o2bb2a_1 _1434_ (.A1_N(_0090_),
    .A2_N(_0077_),
    .B1(_0107_),
    .B2(_0130_),
    .X(_0513_));
 sky130_fd_sc_hd__o21ba_1 _1435_ (.A1(_0416_),
    .A2(_0513_),
    .B1_N(_0445_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _1436_ (.A0(_0486_),
    .A1(_0407_),
    .S(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__or2_1 _1437_ (.A(_0152_),
    .B(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__xor2_1 _1438_ (.A(_0512_),
    .B(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__a31o_1 _1439_ (.A1(_0421_),
    .A2(_0077_),
    .A3(_0090_),
    .B1(_0495_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _1440_ (.A0(net45),
    .A1(_0433_),
    .S(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__xnor2_1 _1441_ (.A(_0517_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__a21o_1 _1442_ (.A1(_0505_),
    .A2(_0506_),
    .B1(_0520_),
    .X(_0521_));
 sky130_fd_sc_hd__nand3_1 _1443_ (.A(_0505_),
    .B(_0506_),
    .C(_0520_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _1444_ (.A(_0521_),
    .B(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__and2_1 _1445_ (.A(_0501_),
    .B(_0502_),
    .X(_0524_));
 sky130_fd_sc_hd__inv_2 _1446_ (.A(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__a311o_1 _1447_ (.A1(_0473_),
    .A2(_0474_),
    .A3(_0468_),
    .B1(_0470_),
    .C1(_0503_),
    .X(_0526_));
 sky130_fd_sc_hd__nand2_1 _1448_ (.A(_0525_),
    .B(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__xnor2_2 _1449_ (.A(_0523_),
    .B(_0527_),
    .Y(net29));
 sky130_fd_sc_hd__inv_2 _1450_ (.A(_0522_),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_1 _1451_ (.A(_0512_),
    .B(_0516_),
    .Y(_0529_));
 sky130_fd_sc_hd__and2_1 _1452_ (.A(_0517_),
    .B(_0519_),
    .X(_0530_));
 sky130_fd_sc_hd__nand2_1 _1453_ (.A(_0344_),
    .B(_0387_),
    .Y(_0531_));
 sky130_fd_sc_hd__and2_1 _1454_ (.A(_0388_),
    .B(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__o21ai_1 _1455_ (.A1(_0398_),
    .A2(_0155_),
    .B1(_0395_),
    .Y(_0533_));
 sky130_fd_sc_hd__a22o_1 _1456_ (.A1(_0287_),
    .A2(_0371_),
    .B1(_0533_),
    .B2(_0421_),
    .X(_0534_));
 sky130_fd_sc_hd__xor2_1 _1457_ (.A(_0532_),
    .B(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__nand2_1 _1458_ (.A(_0022_),
    .B(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__nor2_1 _1459_ (.A(_0416_),
    .B(_0181_),
    .Y(_0537_));
 sky130_fd_sc_hd__o21ai_1 _1460_ (.A1(_0445_),
    .A2(_0537_),
    .B1(_0486_),
    .Y(_0538_));
 sky130_fd_sc_hd__o311a_2 _1461_ (.A1(_0187_),
    .A2(_0445_),
    .A3(_0537_),
    .B1(_0538_),
    .C1(_0241_),
    .X(_0539_));
 sky130_fd_sc_hd__xor2_1 _1462_ (.A(_0536_),
    .B(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__o2bb2a_1 _1463_ (.A1_N(_0112_),
    .A2_N(_0433_),
    .B1(_0495_),
    .B2(_0243_),
    .X(_0541_));
 sky130_fd_sc_hd__xor2_1 _1464_ (.A(_0540_),
    .B(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__o21a_1 _1465_ (.A1(_0529_),
    .A2(_0530_),
    .B1(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__nor3_1 _1466_ (.A(_0529_),
    .B(_0530_),
    .C(_0542_),
    .Y(_0544_));
 sky130_fd_sc_hd__or2_1 _1467_ (.A(_0543_),
    .B(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__a311o_1 _1468_ (.A1(_0525_),
    .A2(_0526_),
    .A3(_0521_),
    .B1(_0528_),
    .C1(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__a31o_1 _1469_ (.A1(_0525_),
    .A2(_0526_),
    .A3(_0521_),
    .B1(_0528_),
    .X(_0547_));
 sky130_fd_sc_hd__nand2_1 _1470_ (.A(_0545_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__and2_1 _1471_ (.A(_0546_),
    .B(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__clkbuf_1 _1472_ (.A(_0549_),
    .X(net18));
 sky130_fd_sc_hd__or2b_1 _1473_ (.A(_0536_),
    .B_N(_0539_),
    .X(_0550_));
 sky130_fd_sc_hd__or2_1 _1474_ (.A(_0540_),
    .B(_0541_),
    .X(_0551_));
 sky130_fd_sc_hd__o211a_1 _1475_ (.A1(_0421_),
    .A2(_0370_),
    .B1(_0156_),
    .C1(_0157_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(_0117_),
    .A1(_0387_),
    .S(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__o21ba_1 _1477_ (.A1(_0237_),
    .A2(_0553_),
    .B1_N(_0484_),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _1478_ (.A(_0541_),
    .B(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _1479_ (.A(_0541_),
    .B(_0554_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _1480_ (.A(_0555_),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__xnor2_1 _1481_ (.A(_0539_),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__a21oi_1 _1482_ (.A1(_0550_),
    .A2(_0551_),
    .B1(_0558_),
    .Y(_0559_));
 sky130_fd_sc_hd__and3_1 _1483_ (.A(_0550_),
    .B(_0551_),
    .C(_0558_),
    .X(_0560_));
 sky130_fd_sc_hd__nor2_2 _1484_ (.A(_0559_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__and2b_1 _1485_ (.A_N(_0543_),
    .B(_0546_),
    .X(_0562_));
 sky130_fd_sc_hd__xnor2_4 _1486_ (.A(_0561_),
    .B(_0562_),
    .Y(net19));
 sky130_fd_sc_hd__inv_2 _1487_ (.A(_0555_),
    .Y(_0563_));
 sky130_fd_sc_hd__o21ai_1 _1488_ (.A1(_0539_),
    .A2(_0563_),
    .B1(_0556_),
    .Y(_0564_));
 sky130_fd_sc_hd__or3_1 _1489_ (.A(_0151_),
    .B(_0532_),
    .C(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__nor2_1 _1490_ (.A(_0543_),
    .B(_0559_),
    .Y(_0566_));
 sky130_fd_sc_hd__a21oi_1 _1491_ (.A1(_0546_),
    .A2(_0566_),
    .B1(_0560_),
    .Y(_0567_));
 sky130_fd_sc_hd__o21a_1 _1492_ (.A1(_0151_),
    .A2(_0532_),
    .B1(_0564_),
    .X(_0568_));
 sky130_fd_sc_hd__a21oi_2 _1493_ (.A1(_0565_),
    .A2(_0567_),
    .B1(_0568_),
    .Y(net20));
 sky130_fd_sc_hd__xnor2_2 _1494_ (.A(_0277_),
    .B(_0276_),
    .Y(net21));
 sky130_fd_sc_hd__clkbuf_4 _1495_ (.A(_0825_),
    .X(_0569_));
 sky130_fd_sc_hd__clkbuf_4 _1496_ (.A(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__buf_4 _1497_ (.A(net31),
    .X(_0571_));
 sky130_fd_sc_hd__buf_4 _1498_ (.A(net30),
    .X(_0572_));
 sky130_fd_sc_hd__xnor2_1 _1499_ (.A(_0571_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__buf_4 _1500_ (.A(net31),
    .X(_0574_));
 sky130_fd_sc_hd__buf_4 _1501_ (.A(_0825_),
    .X(_0575_));
 sky130_fd_sc_hd__nand3_2 _1502_ (.A(_0574_),
    .B(_0572_),
    .C(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__buf_2 _1503_ (.A(net33),
    .X(_0577_));
 sky130_fd_sc_hd__buf_2 _1504_ (.A(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__o211a_1 _1505_ (.A1(_0570_),
    .A2(_0573_),
    .B1(_0576_),
    .C1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__nor2b_2 _1506_ (.A(_0878_),
    .B_N(_0569_),
    .Y(_0580_));
 sky130_fd_sc_hd__nor2_1 _1507_ (.A(_0578_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__or2_1 _1508_ (.A(_0579_),
    .B(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__clkbuf_4 _1509_ (.A(_0577_),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_2 _1510_ (.A(_0572_),
    .B(_0569_),
    .Y(_0584_));
 sky130_fd_sc_hd__or3b_2 _1511_ (.A(_0900_),
    .B(_0825_),
    .C_N(_0878_),
    .X(_0585_));
 sky130_fd_sc_hd__and2_1 _1512_ (.A(_0584_),
    .B(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__buf_2 _1513_ (.A(_0900_),
    .X(_0587_));
 sky130_fd_sc_hd__o21a_2 _1514_ (.A1(_0587_),
    .A2(_0575_),
    .B1(_0577_),
    .X(_0588_));
 sky130_fd_sc_hd__clkbuf_4 _1515_ (.A(net34),
    .X(_0589_));
 sky130_fd_sc_hd__clkbuf_4 _1516_ (.A(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__and2_1 _1517_ (.A(_0571_),
    .B(_0900_),
    .X(_0591_));
 sky130_fd_sc_hd__o21ai_1 _1518_ (.A1(_0587_),
    .A2(_0570_),
    .B1(_0577_),
    .Y(_0592_));
 sky130_fd_sc_hd__or3_1 _1519_ (.A(_0591_),
    .B(_0580_),
    .C(_0592_),
    .X(_0593_));
 sky130_fd_sc_hd__o221ai_2 _1520_ (.A1(_0583_),
    .A2(_0586_),
    .B1(_0588_),
    .B2(_0590_),
    .C1(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__clkbuf_4 _1521_ (.A(_0857_),
    .X(_0595_));
 sky130_fd_sc_hd__a221o_4 _1522_ (.A1(_0868_),
    .A2(_0582_),
    .B1(_0594_),
    .B2(_0595_),
    .C1(_0942_),
    .X(_0596_));
 sky130_fd_sc_hd__clkbuf_2 _1523_ (.A(\p_shaping_I.counter[1] ),
    .X(_0597_));
 sky130_fd_sc_hd__nor2_4 _1524_ (.A(_0571_),
    .B(_0572_),
    .Y(_0598_));
 sky130_fd_sc_hd__buf_2 _1525_ (.A(_0803_),
    .X(_0599_));
 sky130_fd_sc_hd__clkbuf_4 _1526_ (.A(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__nand2_1 _1527_ (.A(_0600_),
    .B(_0868_),
    .Y(_0601_));
 sky130_fd_sc_hd__nand2_1 _1528_ (.A(_0595_),
    .B(_0589_),
    .Y(_0602_));
 sky130_fd_sc_hd__a21oi_4 _1529_ (.A1(_0571_),
    .A2(_0900_),
    .B1(_0569_),
    .Y(_0603_));
 sky130_fd_sc_hd__a21boi_2 _1530_ (.A1(_0878_),
    .A2(_0825_),
    .B1_N(_0900_),
    .Y(_0604_));
 sky130_fd_sc_hd__or2_1 _1531_ (.A(_0803_),
    .B(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__o31a_1 _1532_ (.A1(_0578_),
    .A2(_0598_),
    .A3(_0603_),
    .B1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__inv_2 _1533_ (.A(_0571_),
    .Y(_0607_));
 sky130_fd_sc_hd__inv_2 _1534_ (.A(_0825_),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_1 _1535_ (.A(_0574_),
    .B(_0587_),
    .Y(_0609_));
 sky130_fd_sc_hd__o21a_1 _1536_ (.A1(_0571_),
    .A2(_0900_),
    .B1(_0575_),
    .X(_0610_));
 sky130_fd_sc_hd__a221o_1 _1537_ (.A1(_0607_),
    .A2(_0608_),
    .B1(_0609_),
    .B2(_0610_),
    .C1(_0599_),
    .X(_0611_));
 sky130_fd_sc_hd__nor2b_4 _1538_ (.A(_0575_),
    .B_N(_0572_),
    .Y(_0612_));
 sky130_fd_sc_hd__and2b_2 _1539_ (.A_N(_0825_),
    .B(_0878_),
    .X(_0613_));
 sky130_fd_sc_hd__nor2_2 _1540_ (.A(net35),
    .B(_0589_),
    .Y(_0614_));
 sky130_fd_sc_hd__o31a_1 _1541_ (.A1(_0578_),
    .A2(_0612_),
    .A3(_0613_),
    .B1(_0614_),
    .X(_0615_));
 sky130_fd_sc_hd__nand2_1 _1542_ (.A(_0611_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__o221a_2 _1543_ (.A1(_0598_),
    .A2(_0601_),
    .B1(_0602_),
    .B2(_0606_),
    .C1(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _1544_ (.A(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__or2b_2 _1545_ (.A(_0825_),
    .B_N(_0878_),
    .X(_0619_));
 sky130_fd_sc_hd__nand2b_4 _1546_ (.A_N(_0878_),
    .B(_0569_),
    .Y(_0620_));
 sky130_fd_sc_hd__and3_1 _1547_ (.A(_0600_),
    .B(_0619_),
    .C(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__nor2_1 _1548_ (.A(_0600_),
    .B(_0619_),
    .Y(_0622_));
 sky130_fd_sc_hd__o41a_2 _1549_ (.A1(_0878_),
    .A2(_0900_),
    .A3(_0889_),
    .A4(_0569_),
    .B1(net34),
    .X(_0623_));
 sky130_fd_sc_hd__or2_1 _1550_ (.A(_0595_),
    .B(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__o21bai_1 _1551_ (.A1(_0621_),
    .A2(_0622_),
    .B1_N(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__inv_2 _1552_ (.A(net34),
    .Y(_0626_));
 sky130_fd_sc_hd__clkbuf_4 _1553_ (.A(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__a211o_1 _1554_ (.A1(_0584_),
    .A2(_0585_),
    .B1(_0577_),
    .C1(_0580_),
    .X(_0628_));
 sky130_fd_sc_hd__xor2_4 _1555_ (.A(net31),
    .B(net30),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_4 _1556_ (.A(_0629_),
    .X(_0630_));
 sky130_fd_sc_hd__a21bo_2 _1557_ (.A1(_0571_),
    .A2(_0569_),
    .B1_N(_0889_),
    .X(_0631_));
 sky130_fd_sc_hd__or2_1 _1558_ (.A(_0630_),
    .B(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__a21o_1 _1559_ (.A1(_0571_),
    .A2(_0569_),
    .B1(_0889_),
    .X(_0633_));
 sky130_fd_sc_hd__o221a_1 _1560_ (.A1(_0599_),
    .A2(_0584_),
    .B1(_0633_),
    .B2(_0598_),
    .C1(_0589_),
    .X(_0634_));
 sky130_fd_sc_hd__clkbuf_4 _1561_ (.A(net35),
    .X(_0635_));
 sky130_fd_sc_hd__a311o_1 _1562_ (.A1(_0627_),
    .A2(_0628_),
    .A3(_0632_),
    .B1(_0634_),
    .C1(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__nand2_1 _1563_ (.A(_0625_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__a21oi_1 _1564_ (.A1(_0597_),
    .A2(_0618_),
    .B1(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2_1 _1565_ (.A(\p_shaping_I.counter[1] ),
    .B(\p_shaping_I.counter[0] ),
    .Y(_0639_));
 sky130_fd_sc_hd__buf_2 _1566_ (.A(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__and3_1 _1567_ (.A(_0597_),
    .B(_0637_),
    .C(_0618_),
    .X(_0641_));
 sky130_fd_sc_hd__or3_4 _1568_ (.A(_0638_),
    .B(_0640_),
    .C(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__xor2_4 _1569_ (.A(_0596_),
    .B(_0642_),
    .X(net4));
 sky130_fd_sc_hd__buf_2 _1570_ (.A(\p_shaping_I.bit_in_2 ),
    .X(_0643_));
 sky130_fd_sc_hd__nor2_2 _1571_ (.A(_0635_),
    .B(_0626_),
    .Y(_0644_));
 sky130_fd_sc_hd__and2b_1 _1572_ (.A_N(net31),
    .B(net30),
    .X(_0645_));
 sky130_fd_sc_hd__nand3b_2 _1573_ (.A_N(_0878_),
    .B(_0889_),
    .C(_0569_),
    .Y(_0646_));
 sky130_fd_sc_hd__o32a_1 _1574_ (.A1(_0577_),
    .A2(_0575_),
    .A3(_0645_),
    .B1(_0646_),
    .B2(_0587_),
    .X(_0647_));
 sky130_fd_sc_hd__o21a_1 _1575_ (.A1(_0623_),
    .A2(_0647_),
    .B1(_0635_),
    .X(_0648_));
 sky130_fd_sc_hd__nand2_1 _1576_ (.A(_0620_),
    .B(_0588_),
    .Y(_0649_));
 sky130_fd_sc_hd__a21o_2 _1577_ (.A1(_0570_),
    .A2(_0629_),
    .B1(_0577_),
    .X(_0650_));
 sky130_fd_sc_hd__or2_2 _1578_ (.A(net35),
    .B(_0589_),
    .X(_0651_));
 sky130_fd_sc_hd__a21oi_1 _1579_ (.A1(_0649_),
    .A2(_0650_),
    .B1(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__a311o_2 _1580_ (.A1(_0583_),
    .A2(_0630_),
    .A3(_0644_),
    .B1(_0648_),
    .C1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__and2_1 _1581_ (.A(_0617_),
    .B(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__and2b_1 _1582_ (.A_N(_0889_),
    .B(_0569_),
    .X(_0655_));
 sky130_fd_sc_hd__nand2_2 _1583_ (.A(_0635_),
    .B(_0627_),
    .Y(_0656_));
 sky130_fd_sc_hd__and2b_1 _1584_ (.A_N(_0572_),
    .B(_0571_),
    .X(_0657_));
 sky130_fd_sc_hd__o21a_1 _1585_ (.A1(_0583_),
    .A2(_0657_),
    .B1(_0584_),
    .X(_0658_));
 sky130_fd_sc_hd__o32a_1 _1586_ (.A1(_0577_),
    .A2(_0575_),
    .A3(_0645_),
    .B1(_0603_),
    .B2(_0814_),
    .X(_0659_));
 sky130_fd_sc_hd__clkbuf_4 _1587_ (.A(_0608_),
    .X(_0660_));
 sky130_fd_sc_hd__a31o_1 _1588_ (.A1(_0599_),
    .A2(_0660_),
    .A3(_0591_),
    .B1(_0626_),
    .X(_0661_));
 sky130_fd_sc_hd__and2_1 _1589_ (.A(_0889_),
    .B(_0825_),
    .X(_0662_));
 sky130_fd_sc_hd__nor2_1 _1590_ (.A(_0572_),
    .B(_0575_),
    .Y(_0663_));
 sky130_fd_sc_hd__a2111o_1 _1591_ (.A1(_0645_),
    .A2(_0662_),
    .B1(net34),
    .C1(_0613_),
    .D1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__a21o_2 _1592_ (.A1(_0572_),
    .A2(_0575_),
    .B1(_0889_),
    .X(_0665_));
 sky130_fd_sc_hd__inv_2 _1593_ (.A(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__o22a_1 _1594_ (.A1(_0659_),
    .A2(_0661_),
    .B1(_0664_),
    .B2(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_4 _1595_ (.A(_0635_),
    .X(_0668_));
 sky130_fd_sc_hd__o32a_1 _1596_ (.A1(_0655_),
    .A2(_0656_),
    .A3(_0658_),
    .B1(_0667_),
    .B2(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__or3_1 _1597_ (.A(_0643_),
    .B(_0654_),
    .C(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__o21ai_1 _1598_ (.A1(_0643_),
    .A2(_0654_),
    .B1(_0669_),
    .Y(_0671_));
 sky130_fd_sc_hd__o21ai_1 _1599_ (.A1(_0583_),
    .A2(_0932_),
    .B1(_0590_),
    .Y(_0672_));
 sky130_fd_sc_hd__nor2_4 _1600_ (.A(_0575_),
    .B(_0629_),
    .Y(_0673_));
 sky130_fd_sc_hd__or2b_1 _1601_ (.A(_0878_),
    .B_N(_0900_),
    .X(_0674_));
 sky130_fd_sc_hd__nor2_1 _1602_ (.A(_0660_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__a2111o_1 _1603_ (.A1(_0578_),
    .A2(_0610_),
    .B1(_0673_),
    .C1(_0675_),
    .D1(_0589_),
    .X(_0676_));
 sky130_fd_sc_hd__nor2_1 _1604_ (.A(_0574_),
    .B(_0578_),
    .Y(_0677_));
 sky130_fd_sc_hd__a21o_1 _1605_ (.A1(_0578_),
    .A2(_0576_),
    .B1(net35),
    .X(_0678_));
 sky130_fd_sc_hd__o31ai_1 _1606_ (.A1(_0677_),
    .A2(_0655_),
    .A3(_0678_),
    .B1(_0651_),
    .Y(_0679_));
 sky130_fd_sc_hd__inv_2 _1607_ (.A(_0572_),
    .Y(_0680_));
 sky130_fd_sc_hd__a31o_1 _1608_ (.A1(_0680_),
    .A2(_0619_),
    .A3(_0620_),
    .B1(_0578_),
    .X(_0681_));
 sky130_fd_sc_hd__nand3_1 _1609_ (.A(_0627_),
    .B(_0586_),
    .C(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__a32o_1 _1610_ (.A1(_0668_),
    .A2(_0672_),
    .A3(_0676_),
    .B1(_0679_),
    .B2(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__inv_2 _1611_ (.A(\p_shaping_I.bit_in_1 ),
    .Y(_0684_));
 sky130_fd_sc_hd__o21a_1 _1612_ (.A1(_0637_),
    .A2(_0683_),
    .B1(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__o31a_1 _1613_ (.A1(_0599_),
    .A2(_0580_),
    .A3(_0645_),
    .B1(_0626_),
    .X(_0686_));
 sky130_fd_sc_hd__a21o_1 _1614_ (.A1(_0589_),
    .A2(_0910_),
    .B1(_0595_),
    .X(_0687_));
 sky130_fd_sc_hd__a21o_1 _1615_ (.A1(_0650_),
    .A2(_0686_),
    .B1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__a211o_1 _1616_ (.A1(_0570_),
    .A2(_0629_),
    .B1(_0663_),
    .C1(_0577_),
    .X(_0689_));
 sky130_fd_sc_hd__a2bb2o_1 _1617_ (.A1_N(_0587_),
    .A2_N(_0631_),
    .B1(_0657_),
    .B2(_0655_),
    .X(_0690_));
 sky130_fd_sc_hd__a221o_1 _1618_ (.A1(_0686_),
    .A2(_0689_),
    .B1(_0690_),
    .B2(_0589_),
    .C1(_0635_),
    .X(_0691_));
 sky130_fd_sc_hd__nand2_1 _1619_ (.A(_0688_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _1620_ (.A(\p_shaping_I.ctl_1 ),
    .B(net48),
    .Y(_0693_));
 sky130_fd_sc_hd__xnor2_1 _1621_ (.A(\p_shaping_I.bit_in ),
    .B(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__nand2_2 _1622_ (.A(net42),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_1 _1623_ (.A(_0692_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__xnor2_1 _1624_ (.A(_0685_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__a31oi_1 _1625_ (.A1(_0597_),
    .A2(_0670_),
    .A3(_0671_),
    .B1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__and4_1 _1626_ (.A(_0597_),
    .B(_0670_),
    .C(_0671_),
    .D(_0697_),
    .X(_0699_));
 sky130_fd_sc_hd__clkbuf_4 _1627_ (.A(_0590_),
    .X(_0700_));
 sky130_fd_sc_hd__o31a_1 _1628_ (.A1(_0680_),
    .A2(_0583_),
    .A3(_0613_),
    .B1(_0635_),
    .X(_0701_));
 sky130_fd_sc_hd__buf_2 _1629_ (.A(_0583_),
    .X(_0702_));
 sky130_fd_sc_hd__a21oi_1 _1630_ (.A1(_0932_),
    .A2(_0604_),
    .B1(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__o2bb2a_1 _1631_ (.A1_N(_0605_),
    .A2_N(_0701_),
    .B1(_0703_),
    .B2(_0678_),
    .X(_0704_));
 sky130_fd_sc_hd__nand2b_1 _1632_ (.A_N(_0572_),
    .B(_0575_),
    .Y(_0705_));
 sky130_fd_sc_hd__and2_2 _1633_ (.A(_0578_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__a211o_1 _1634_ (.A1(_0620_),
    .A2(_0706_),
    .B1(_0673_),
    .C1(_0602_),
    .X(_0707_));
 sky130_fd_sc_hd__o21ai_1 _1635_ (.A1(_0700_),
    .A2(_0704_),
    .B1(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__o211ai_1 _1636_ (.A1(_0603_),
    .A2(_0650_),
    .B1(_0868_),
    .C1(_0649_),
    .Y(_0709_));
 sky130_fd_sc_hd__or2b_1 _1637_ (.A(_0900_),
    .B_N(_0571_),
    .X(_0710_));
 sky130_fd_sc_hd__mux2_1 _1638_ (.A0(_0576_),
    .A1(_0710_),
    .S(_0599_),
    .X(_0711_));
 sky130_fd_sc_hd__or3_1 _1639_ (.A(_0635_),
    .B(_0590_),
    .C(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__and2_1 _1640_ (.A(_0583_),
    .B(_0932_),
    .X(_0713_));
 sky130_fd_sc_hd__and3_1 _1641_ (.A(_0599_),
    .B(_0620_),
    .C(_0674_),
    .X(_0714_));
 sky130_fd_sc_hd__o21ai_1 _1642_ (.A1(_0713_),
    .A2(_0714_),
    .B1(_0644_),
    .Y(_0715_));
 sky130_fd_sc_hd__and3_2 _1643_ (.A(_0709_),
    .B(_0712_),
    .C(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__a21oi_1 _1644_ (.A1(_0596_),
    .A2(_0716_),
    .B1(\p_shaping_I.bit_in ),
    .Y(_0717_));
 sky130_fd_sc_hd__xnor2_1 _1645_ (.A(_0708_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__or4_1 _1646_ (.A(_0640_),
    .B(_0698_),
    .C(_0699_),
    .D(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__o31ai_1 _1647_ (.A1(_0640_),
    .A2(_0698_),
    .A3(_0699_),
    .B1(_0718_),
    .Y(_0720_));
 sky130_fd_sc_hd__clkinv_2 _1648_ (.A(_0639_),
    .Y(_0025_));
 sky130_fd_sc_hd__o21ai_1 _1649_ (.A1(_0643_),
    .A2(_0617_),
    .B1(_0653_),
    .Y(_0721_));
 sky130_fd_sc_hd__or3_1 _1650_ (.A(\p_shaping_I.bit_in_2 ),
    .B(_0617_),
    .C(_0653_),
    .X(_0722_));
 sky130_fd_sc_hd__a21o_1 _1651_ (.A1(_0625_),
    .A2(_0636_),
    .B1(\p_shaping_I.bit_in_1 ),
    .X(_0723_));
 sky130_fd_sc_hd__xnor2_1 _1652_ (.A(_0723_),
    .B(_0683_),
    .Y(_0724_));
 sky130_fd_sc_hd__nand4_1 _1653_ (.A(_0597_),
    .B(_0721_),
    .C(_0722_),
    .D(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__a31o_1 _1654_ (.A1(_0597_),
    .A2(_0721_),
    .A3(_0722_),
    .B1(_0724_),
    .X(_0726_));
 sky130_fd_sc_hd__and3_1 _1655_ (.A(_0025_),
    .B(_0725_),
    .C(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__nor2_1 _1656_ (.A(_0114_),
    .B(_0596_),
    .Y(_0728_));
 sky130_fd_sc_hd__xnor2_2 _1657_ (.A(_0716_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__a21bo_1 _1658_ (.A1(_0727_),
    .A2(_0729_),
    .B1_N(_0725_),
    .X(_0730_));
 sky130_fd_sc_hd__a21o_1 _1659_ (.A1(_0719_),
    .A2(_0720_),
    .B1(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__and3_1 _1660_ (.A(_0719_),
    .B(_0720_),
    .C(_0730_),
    .X(_0732_));
 sky130_fd_sc_hd__inv_2 _1661_ (.A(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_2 _1662_ (.A(_0731_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__xnor2_2 _1663_ (.A(_0727_),
    .B(_0729_),
    .Y(_0735_));
 sky130_fd_sc_hd__o21bai_4 _1664_ (.A1(_0596_),
    .A2(_0642_),
    .B1_N(_0641_),
    .Y(_0736_));
 sky130_fd_sc_hd__and2b_1 _1665_ (.A_N(_0735_),
    .B(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__xnor2_4 _1666_ (.A(_0734_),
    .B(_0737_),
    .Y(net9));
 sky130_fd_sc_hd__and3_1 _1667_ (.A(_0617_),
    .B(_0653_),
    .C(_0669_),
    .X(_0738_));
 sky130_fd_sc_hd__a211o_1 _1668_ (.A1(_0570_),
    .A2(_0710_),
    .B1(_0613_),
    .C1(_0599_),
    .X(_0739_));
 sky130_fd_sc_hd__a311o_1 _1669_ (.A1(_0619_),
    .A2(_0620_),
    .A3(_0584_),
    .B1(_0598_),
    .C1(_0577_),
    .X(_0740_));
 sky130_fd_sc_hd__o211ai_1 _1670_ (.A1(_0814_),
    .A2(_0603_),
    .B1(_0588_),
    .C1(_0620_),
    .Y(_0741_));
 sky130_fd_sc_hd__o21a_1 _1671_ (.A1(_0612_),
    .A2(_0633_),
    .B1(_0626_),
    .X(_0742_));
 sky130_fd_sc_hd__a32o_1 _1672_ (.A1(_0589_),
    .A2(_0739_),
    .A3(_0740_),
    .B1(_0741_),
    .B2(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__a21oi_1 _1673_ (.A1(_0570_),
    .A2(_0630_),
    .B1(_0612_),
    .Y(_0744_));
 sky130_fd_sc_hd__xor2_1 _1674_ (.A(_0714_),
    .B(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__o2bb2a_1 _1675_ (.A1_N(_0595_),
    .A2_N(_0743_),
    .B1(_0745_),
    .B2(_0656_),
    .X(_0746_));
 sky130_fd_sc_hd__o21ai_1 _1676_ (.A1(_0643_),
    .A2(_0738_),
    .B1(_0746_),
    .Y(_0747_));
 sky130_fd_sc_hd__or3_1 _1677_ (.A(_0643_),
    .B(_0746_),
    .C(_0738_),
    .X(_0748_));
 sky130_fd_sc_hd__o31a_1 _1678_ (.A1(_0637_),
    .A2(_0683_),
    .A3(_0692_),
    .B1(_0684_),
    .X(_0749_));
 sky130_fd_sc_hd__and2_1 _1679_ (.A(net42),
    .B(_0694_),
    .X(_0750_));
 sky130_fd_sc_hd__clkbuf_2 _1680_ (.A(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__a21o_1 _1681_ (.A1(_0660_),
    .A2(_0573_),
    .B1(_0610_),
    .X(_0752_));
 sky130_fd_sc_hd__a21oi_1 _1682_ (.A1(_0702_),
    .A2(_0752_),
    .B1(_0581_),
    .Y(_0753_));
 sky130_fd_sc_hd__a31o_1 _1683_ (.A1(_0619_),
    .A2(_0620_),
    .A3(_0584_),
    .B1(_0578_),
    .X(_0754_));
 sky130_fd_sc_hd__and3_1 _1684_ (.A(_0627_),
    .B(_0611_),
    .C(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__a31o_1 _1685_ (.A1(_0590_),
    .A2(_0605_),
    .A3(_0665_),
    .B1(_0635_),
    .X(_0756_));
 sky130_fd_sc_hd__o22ai_2 _1686_ (.A1(_0624_),
    .A2(_0753_),
    .B1(_0755_),
    .B2(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__nor2_1 _1687_ (.A(_0751_),
    .B(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__xnor2_1 _1688_ (.A(_0749_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__a31oi_1 _1689_ (.A1(_0597_),
    .A2(_0747_),
    .A3(_0748_),
    .B1(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__and4_1 _1690_ (.A(_0597_),
    .B(_0747_),
    .C(_0748_),
    .D(_0759_),
    .X(_0761_));
 sky130_fd_sc_hd__or3_1 _1691_ (.A(_0640_),
    .B(_0760_),
    .C(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__nor2_1 _1692_ (.A(_0627_),
    .B(_0910_),
    .Y(_0763_));
 sky130_fd_sc_hd__a221oi_1 _1693_ (.A1(_0630_),
    .A2(_0588_),
    .B1(_0673_),
    .B2(_0600_),
    .C1(_0700_),
    .Y(_0764_));
 sky130_fd_sc_hd__o21a_1 _1694_ (.A1(_0763_),
    .A2(_0764_),
    .B1(_0668_),
    .X(_0765_));
 sky130_fd_sc_hd__nand2_2 _1695_ (.A(_0660_),
    .B(_0598_),
    .Y(_0766_));
 sky130_fd_sc_hd__o221a_1 _1696_ (.A1(_0587_),
    .A2(_0646_),
    .B1(_0706_),
    .B2(_0598_),
    .C1(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__nor2_1 _1697_ (.A(_0660_),
    .B(_0657_),
    .Y(_0768_));
 sky130_fd_sc_hd__o211a_1 _1698_ (.A1(_0702_),
    .A2(_0768_),
    .B1(_0605_),
    .C1(_0595_),
    .X(_0769_));
 sky130_fd_sc_hd__o2bb2a_1 _1699_ (.A1_N(_0700_),
    .A2_N(_0767_),
    .B1(_0769_),
    .B2(_0644_),
    .X(_0770_));
 sky130_fd_sc_hd__nor2_2 _1700_ (.A(_0765_),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__and3b_1 _1701_ (.A_N(_0708_),
    .B(_0716_),
    .C(_0596_),
    .X(_0772_));
 sky130_fd_sc_hd__or2_1 _1702_ (.A(_0114_),
    .B(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__xnor2_1 _1703_ (.A(_0771_),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__xnor2_1 _1704_ (.A(_0762_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__or2b_1 _1705_ (.A(_0699_),
    .B_N(_0719_),
    .X(_0776_));
 sky130_fd_sc_hd__and2b_1 _1706_ (.A_N(_0775_),
    .B(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__or2b_1 _1707_ (.A(_0776_),
    .B_N(_0775_),
    .X(_0778_));
 sky130_fd_sc_hd__and2b_1 _1708_ (.A_N(_0777_),
    .B(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__a21o_2 _1709_ (.A1(_0731_),
    .A2(_0737_),
    .B1(_0732_),
    .X(_0780_));
 sky130_fd_sc_hd__xor2_2 _1710_ (.A(_0779_),
    .B(_0780_),
    .X(net10));
 sky130_fd_sc_hd__buf_2 _1711_ (.A(_0597_),
    .X(_0781_));
 sky130_fd_sc_hd__a41o_1 _1712_ (.A1(_0617_),
    .A2(_0653_),
    .A3(_0669_),
    .A4(_0746_),
    .B1(\p_shaping_I.bit_in_2 ),
    .X(_0782_));
 sky130_fd_sc_hd__a21oi_2 _1713_ (.A1(_0574_),
    .A2(_0570_),
    .B1(_0583_),
    .Y(_0783_));
 sky130_fd_sc_hd__a21o_1 _1714_ (.A1(_0583_),
    .A2(_0609_),
    .B1(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__o211a_1 _1715_ (.A1(_0630_),
    .A2(_0631_),
    .B1(_0650_),
    .C1(_0635_),
    .X(_0785_));
 sky130_fd_sc_hd__o211ai_1 _1716_ (.A1(_0607_),
    .A2(_0612_),
    .B1(_0705_),
    .C1(_0583_),
    .Y(_0786_));
 sky130_fd_sc_hd__a31oi_1 _1717_ (.A1(_0595_),
    .A2(_0689_),
    .A3(_0786_),
    .B1(_0627_),
    .Y(_0787_));
 sky130_fd_sc_hd__a211o_1 _1718_ (.A1(_0614_),
    .A2(_0784_),
    .B1(_0785_),
    .C1(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__xor2_1 _1719_ (.A(_0782_),
    .B(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__and2_1 _1720_ (.A(_0684_),
    .B(_0757_),
    .X(_0790_));
 sky130_fd_sc_hd__nand2_1 _1721_ (.A(_0570_),
    .B(_0630_),
    .Y(_0791_));
 sky130_fd_sc_hd__nand2_1 _1722_ (.A(_0588_),
    .B(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__or2_1 _1723_ (.A(_0660_),
    .B(_0598_),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_1 _1724_ (.A(_0932_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hd__a31o_1 _1725_ (.A1(_0627_),
    .A2(_0792_),
    .A3(_0794_),
    .B1(_0623_),
    .X(_0795_));
 sky130_fd_sc_hd__or4_1 _1726_ (.A(_0590_),
    .B(_0677_),
    .C(_0580_),
    .D(_0622_),
    .X(_0796_));
 sky130_fd_sc_hd__o211a_1 _1727_ (.A1(_0702_),
    .A2(_0585_),
    .B1(_0674_),
    .C1(_0590_),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_1 _1728_ (.A(_0668_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__a22o_1 _1729_ (.A1(_0668_),
    .A2(_0795_),
    .B1(_0796_),
    .B2(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__o21bai_1 _1730_ (.A1(_0749_),
    .A2(_0790_),
    .B1_N(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__or3b_1 _1731_ (.A(_0749_),
    .B(_0790_),
    .C_N(_0799_),
    .X(_0801_));
 sky130_fd_sc_hd__a21oi_1 _1732_ (.A1(_0592_),
    .A2(_0681_),
    .B1(_0656_),
    .Y(_0802_));
 sky130_fd_sc_hd__o211a_1 _1733_ (.A1(_0660_),
    .A2(_0674_),
    .B1(_0710_),
    .C1(_0599_),
    .X(_0804_));
 sky130_fd_sc_hd__a2bb2o_1 _1734_ (.A1_N(_0587_),
    .A2_N(_0631_),
    .B1(_0603_),
    .B2(_0599_),
    .X(_0805_));
 sky130_fd_sc_hd__o211a_1 _1735_ (.A1(_0706_),
    .A2(_0804_),
    .B1(_0805_),
    .C1(_0644_),
    .X(_0806_));
 sky130_fd_sc_hd__nor2_1 _1736_ (.A(_0651_),
    .B(_0805_),
    .Y(_0807_));
 sky130_fd_sc_hd__or3_1 _1737_ (.A(_0802_),
    .B(_0806_),
    .C(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__o31a_2 _1738_ (.A1(_0692_),
    .A2(_0757_),
    .A3(_0808_),
    .B1(_0684_),
    .X(_0809_));
 sky130_fd_sc_hd__nor2_1 _1739_ (.A(_0695_),
    .B(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__a31o_1 _1740_ (.A1(_0695_),
    .A2(_0800_),
    .A3(_0801_),
    .B1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__a21oi_1 _1741_ (.A1(_0781_),
    .A2(_0789_),
    .B1(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__and3_1 _1742_ (.A(_0781_),
    .B(_0789_),
    .C(_0811_),
    .X(_0813_));
 sky130_fd_sc_hd__o311a_1 _1743_ (.A1(_0574_),
    .A2(_0600_),
    .A3(_0612_),
    .B1(_0665_),
    .C1(_0700_),
    .X(_0815_));
 sky130_fd_sc_hd__a21oi_1 _1744_ (.A1(_0574_),
    .A2(_0633_),
    .B1(_0700_),
    .Y(_0816_));
 sky130_fd_sc_hd__clkbuf_4 _1745_ (.A(_0702_),
    .X(_0817_));
 sky130_fd_sc_hd__or2_1 _1746_ (.A(_0603_),
    .B(_0610_),
    .X(_0818_));
 sky130_fd_sc_hd__or2_1 _1747_ (.A(_0587_),
    .B(_0570_),
    .X(_0819_));
 sky130_fd_sc_hd__and3_1 _1748_ (.A(_0600_),
    .B(_0609_),
    .C(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__a21o_1 _1749_ (.A1(_0817_),
    .A2(_0818_),
    .B1(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__o32a_1 _1750_ (.A1(_0668_),
    .A2(_0815_),
    .A3(_0816_),
    .B1(_0821_),
    .B2(_0656_),
    .X(_0822_));
 sky130_fd_sc_hd__a21o_1 _1751_ (.A1(_0771_),
    .A2(_0772_),
    .B1(_0114_),
    .X(_0823_));
 sky130_fd_sc_hd__xnor2_1 _1752_ (.A(_0822_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__or4_2 _1753_ (.A(_0640_),
    .B(_0812_),
    .C(_0813_),
    .D(_0824_),
    .X(_0826_));
 sky130_fd_sc_hd__o31ai_2 _1754_ (.A1(_0640_),
    .A2(_0812_),
    .A3(_0813_),
    .B1(_0824_),
    .Y(_0827_));
 sky130_fd_sc_hd__o21bai_2 _1755_ (.A1(_0762_),
    .A2(_0774_),
    .B1_N(_0761_),
    .Y(_0828_));
 sky130_fd_sc_hd__nand3_4 _1756_ (.A(_0826_),
    .B(_0827_),
    .C(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__a21o_1 _1757_ (.A1(_0826_),
    .A2(_0827_),
    .B1(_0828_),
    .X(_0830_));
 sky130_fd_sc_hd__o2111ai_4 _1758_ (.A1(_0777_),
    .A2(_0780_),
    .B1(_0829_),
    .C1(_0830_),
    .D1(_0778_),
    .Y(_0831_));
 sky130_fd_sc_hd__or2_1 _1759_ (.A(_0777_),
    .B(_0780_),
    .X(_0832_));
 sky130_fd_sc_hd__a22o_1 _1760_ (.A1(_0829_),
    .A2(_0830_),
    .B1(_0832_),
    .B2(_0778_),
    .X(_0833_));
 sky130_fd_sc_hd__and2_1 _1761_ (.A(_0831_),
    .B(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_1 _1762_ (.A(_0834_),
    .X(net11));
 sky130_fd_sc_hd__inv_2 _1763_ (.A(_0813_),
    .Y(_0836_));
 sky130_fd_sc_hd__or2_1 _1764_ (.A(\p_shaping_I.bit_in_2 ),
    .B(_0788_),
    .X(_0837_));
 sky130_fd_sc_hd__inv_2 _1765_ (.A(_0706_),
    .Y(_0838_));
 sky130_fd_sc_hd__or3b_1 _1766_ (.A(_0633_),
    .B(_0598_),
    .C_N(_0932_),
    .X(_0839_));
 sky130_fd_sc_hd__o211a_1 _1767_ (.A1(_0630_),
    .A2(_0631_),
    .B1(_0839_),
    .C1(_0590_),
    .X(_0840_));
 sky130_fd_sc_hd__or2_1 _1768_ (.A(_0600_),
    .B(_0603_),
    .X(_0841_));
 sky130_fd_sc_hd__o21ai_1 _1769_ (.A1(_0702_),
    .A2(_0814_),
    .B1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__o21a_1 _1770_ (.A1(_0590_),
    .A2(_0842_),
    .B1(_0668_),
    .X(_0843_));
 sky130_fd_sc_hd__a311o_1 _1771_ (.A1(_0628_),
    .A2(_0614_),
    .A3(_0838_),
    .B1(_0840_),
    .C1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__a21o_1 _1772_ (.A1(_0782_),
    .A2(_0837_),
    .B1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__nand3_1 _1773_ (.A(_0782_),
    .B(_0844_),
    .C(_0837_),
    .Y(_0847_));
 sky130_fd_sc_hd__and3_1 _1774_ (.A(_0597_),
    .B(_0845_),
    .C(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__a211oi_1 _1775_ (.A1(_0684_),
    .A2(_0692_),
    .B1(_0808_),
    .C1(_0790_),
    .Y(_0849_));
 sky130_fd_sc_hd__a211oi_1 _1776_ (.A1(_0684_),
    .A2(_0808_),
    .B1(_0849_),
    .C1(_0751_),
    .Y(_0850_));
 sky130_fd_sc_hd__nor3_1 _1777_ (.A(_0810_),
    .B(_0848_),
    .C(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__o21a_1 _1778_ (.A1(_0810_),
    .A2(_0850_),
    .B1(_0848_),
    .X(_0852_));
 sky130_fd_sc_hd__or3_1 _1779_ (.A(_0640_),
    .B(_0851_),
    .C(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__and3_1 _1780_ (.A(_0771_),
    .B(_0772_),
    .C(_0822_),
    .X(_0854_));
 sky130_fd_sc_hd__or2_1 _1781_ (.A(_0114_),
    .B(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__nor2_1 _1782_ (.A(_0700_),
    .B(_0662_),
    .Y(_0856_));
 sky130_fd_sc_hd__o21a_1 _1783_ (.A1(_0665_),
    .A2(_0673_),
    .B1(_0856_),
    .X(_0858_));
 sky130_fd_sc_hd__a21oi_1 _1784_ (.A1(_0677_),
    .A2(_0663_),
    .B1(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__clkbuf_4 _1785_ (.A(_0700_),
    .X(_0860_));
 sky130_fd_sc_hd__a31o_1 _1786_ (.A1(_0817_),
    .A2(_0584_),
    .A3(_0585_),
    .B1(_0783_),
    .X(_0861_));
 sky130_fd_sc_hd__nor2_1 _1787_ (.A(_0860_),
    .B(_0835_),
    .Y(_0862_));
 sky130_fd_sc_hd__a211o_1 _1788_ (.A1(_0860_),
    .A2(_0861_),
    .B1(_0862_),
    .C1(_0668_),
    .X(_0863_));
 sky130_fd_sc_hd__o21a_1 _1789_ (.A1(_0595_),
    .A2(_0859_),
    .B1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__xnor2_1 _1790_ (.A(_0855_),
    .B(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__xnor2_1 _1791_ (.A(_0853_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__a21oi_1 _1792_ (.A1(_0836_),
    .A2(_0826_),
    .B1(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__and3_1 _1793_ (.A(_0836_),
    .B(_0826_),
    .C(_0866_),
    .X(_0869_));
 sky130_fd_sc_hd__or2_1 _1794_ (.A(_0867_),
    .B(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__nand2_1 _1795_ (.A(_0829_),
    .B(_0831_),
    .Y(_0871_));
 sky130_fd_sc_hd__xnor2_1 _1796_ (.A(_0870_),
    .B(_0871_),
    .Y(net12));
 sky130_fd_sc_hd__a21o_1 _1797_ (.A1(_0836_),
    .A2(_0826_),
    .B1(_0866_),
    .X(_0872_));
 sky130_fd_sc_hd__a21o_1 _1798_ (.A1(_0660_),
    .A2(_0591_),
    .B1(_0665_),
    .X(_0873_));
 sky130_fd_sc_hd__o21ai_1 _1799_ (.A1(_0700_),
    .A2(_0646_),
    .B1(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__and3_1 _1800_ (.A(_0590_),
    .B(_0766_),
    .C(_0793_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _1801_ (.A0(_0874_),
    .A1(_0873_),
    .S(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__clkbuf_4 _1802_ (.A(_0668_),
    .X(_0877_));
 sky130_fd_sc_hd__o32a_1 _1803_ (.A1(_0817_),
    .A2(_0814_),
    .A3(_0656_),
    .B1(_0876_),
    .B2(_0877_),
    .X(_0879_));
 sky130_fd_sc_hd__a31o_2 _1804_ (.A1(_0782_),
    .A2(_0788_),
    .A3(_0844_),
    .B1(_0643_),
    .X(_0880_));
 sky130_fd_sc_hd__xor2_1 _1805_ (.A(_0879_),
    .B(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__xnor2_1 _1806_ (.A(_0579_),
    .B(_0604_),
    .Y(_0882_));
 sky130_fd_sc_hd__and4_1 _1807_ (.A(_0607_),
    .B(_0589_),
    .C(_0584_),
    .D(_0819_),
    .X(_0883_));
 sky130_fd_sc_hd__o21ai_1 _1808_ (.A1(_0817_),
    .A2(_0705_),
    .B1(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__or3_1 _1809_ (.A(_0702_),
    .B(_0705_),
    .C(_0883_),
    .X(_0885_));
 sky130_fd_sc_hd__o311a_1 _1810_ (.A1(_0700_),
    .A2(_0673_),
    .A3(_0838_),
    .B1(_0884_),
    .C1(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__o221a_1 _1811_ (.A1(_0656_),
    .A2(_0882_),
    .B1(_0886_),
    .B2(_0877_),
    .C1(_0695_),
    .X(_0887_));
 sky130_fd_sc_hd__xnor2_1 _1812_ (.A(_0809_),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__a21oi_1 _1813_ (.A1(_0781_),
    .A2(_0881_),
    .B1(_0888_),
    .Y(_0890_));
 sky130_fd_sc_hd__and3_1 _1814_ (.A(_0781_),
    .B(_0881_),
    .C(_0888_),
    .X(_0891_));
 sky130_fd_sc_hd__or3_1 _1815_ (.A(_0640_),
    .B(_0890_),
    .C(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__and2_1 _1816_ (.A(_0854_),
    .B(_0864_),
    .X(_0893_));
 sky130_fd_sc_hd__nor2_2 _1817_ (.A(_0114_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__a2111oi_1 _1818_ (.A1(_0630_),
    .A2(_0662_),
    .B1(_0622_),
    .C1(_0627_),
    .D1(_0783_),
    .Y(_0895_));
 sky130_fd_sc_hd__nor2_1 _1819_ (.A(_0706_),
    .B(_0804_),
    .Y(_0896_));
 sky130_fd_sc_hd__o32a_1 _1820_ (.A1(_0877_),
    .A2(_0856_),
    .A3(_0895_),
    .B1(_0656_),
    .B2(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__xnor2_2 _1821_ (.A(_0894_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__xnor2_2 _1822_ (.A(_0892_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__o21bai_2 _1823_ (.A1(_0853_),
    .A2(_0865_),
    .B1_N(_0852_),
    .Y(_0901_));
 sky130_fd_sc_hd__xnor2_2 _1824_ (.A(_0899_),
    .B(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__a311oi_4 _1825_ (.A1(_0829_),
    .A2(_0831_),
    .A3(_0872_),
    .B1(_0869_),
    .C1(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__a31o_1 _1826_ (.A1(_0829_),
    .A2(_0831_),
    .A3(_0872_),
    .B1(_0869_),
    .X(_0904_));
 sky130_fd_sc_hd__nand2_1 _1827_ (.A(_0902_),
    .B(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__and2b_1 _1828_ (.A_N(_0903_),
    .B(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__clkbuf_1 _1829_ (.A(_0906_),
    .X(net13));
 sky130_fd_sc_hd__a21o_1 _1830_ (.A1(_0660_),
    .A2(_0591_),
    .B1(_0580_),
    .X(_0907_));
 sky130_fd_sc_hd__a31o_1 _1831_ (.A1(_0817_),
    .A2(_0860_),
    .A3(_0766_),
    .B1(_0877_),
    .X(_0908_));
 sky130_fd_sc_hd__and2_1 _1832_ (.A(_0689_),
    .B(_0862_),
    .X(_0909_));
 sky130_fd_sc_hd__a211o_1 _1833_ (.A1(_0860_),
    .A2(_0907_),
    .B1(_0908_),
    .C1(_0909_),
    .X(_0911_));
 sky130_fd_sc_hd__nand2_1 _1834_ (.A(_0880_),
    .B(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__or2_1 _1835_ (.A(_0880_),
    .B(_0911_),
    .X(_0913_));
 sky130_fd_sc_hd__or2_1 _1836_ (.A(_0574_),
    .B(_0702_),
    .X(_0914_));
 sky130_fd_sc_hd__a21o_1 _1837_ (.A1(_0914_),
    .A2(_0611_),
    .B1(_0687_),
    .X(_0915_));
 sky130_fd_sc_hd__nor2_1 _1838_ (.A(_0612_),
    .B(_0633_),
    .Y(_0916_));
 sky130_fd_sc_hd__and3_1 _1839_ (.A(_0702_),
    .B(_0766_),
    .C(_0791_),
    .X(_0917_));
 sky130_fd_sc_hd__nand2_1 _1840_ (.A(_0702_),
    .B(_0644_),
    .Y(_0918_));
 sky130_fd_sc_hd__o32a_1 _1841_ (.A1(_0651_),
    .A2(_0916_),
    .A3(_0917_),
    .B1(_0918_),
    .B2(_0768_),
    .X(_0919_));
 sky130_fd_sc_hd__o311a_1 _1842_ (.A1(_0602_),
    .A2(_0650_),
    .A3(_0673_),
    .B1(_0915_),
    .C1(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _1843_ (.A0(\p_shaping_I.bit_in_1 ),
    .A1(_0809_),
    .S(_0920_),
    .X(_0922_));
 sky130_fd_sc_hd__xnor2_1 _1844_ (.A(_0695_),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__a31o_1 _1845_ (.A1(_0781_),
    .A2(_0912_),
    .A3(_0913_),
    .B1(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__nand4_2 _1846_ (.A(_0781_),
    .B(_0923_),
    .C(_0912_),
    .D(_0913_),
    .Y(_0925_));
 sky130_fd_sc_hd__and3_1 _1847_ (.A(_0025_),
    .B(_0924_),
    .C(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__o311a_1 _1848_ (.A1(_0817_),
    .A2(_0814_),
    .A3(_0603_),
    .B1(_0646_),
    .C1(_0627_),
    .X(_0927_));
 sky130_fd_sc_hd__nor2_1 _1849_ (.A(_0763_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__o22a_1 _1850_ (.A1(_0918_),
    .A2(_0794_),
    .B1(_0928_),
    .B2(_0595_),
    .X(_0929_));
 sky130_fd_sc_hd__xor2_2 _1851_ (.A(_0894_),
    .B(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__xnor2_1 _1852_ (.A(_0926_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__nor2_1 _1853_ (.A(_0640_),
    .B(_0890_),
    .Y(_0933_));
 sky130_fd_sc_hd__a21o_1 _1854_ (.A1(_0933_),
    .A2(_0898_),
    .B1(_0891_),
    .X(_0934_));
 sky130_fd_sc_hd__and2_1 _1855_ (.A(_0931_),
    .B(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__nor2_1 _1856_ (.A(_0931_),
    .B(_0934_),
    .Y(_0936_));
 sky130_fd_sc_hd__nor2_2 _1857_ (.A(_0935_),
    .B(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _1858_ (.A(_0899_),
    .B(_0901_),
    .Y(_0938_));
 sky130_fd_sc_hd__inv_2 _1859_ (.A(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__nor2_2 _1860_ (.A(_0939_),
    .B(_0903_),
    .Y(_0940_));
 sky130_fd_sc_hd__xnor2_4 _1861_ (.A(_0937_),
    .B(_0940_),
    .Y(net14));
 sky130_fd_sc_hd__nor2_1 _1862_ (.A(_0650_),
    .B(_0673_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21a_1 _1863_ (.A1(_0623_),
    .A2(_0941_),
    .B1(_0668_),
    .X(_0943_));
 sky130_fd_sc_hd__o311a_1 _1864_ (.A1(_0817_),
    .A2(_0612_),
    .A3(_0598_),
    .B1(_0631_),
    .C1(_0644_),
    .X(_0944_));
 sky130_fd_sc_hd__or3_1 _1865_ (.A(_0700_),
    .B(_0592_),
    .C(_0768_),
    .X(_0945_));
 sky130_fd_sc_hd__o31a_1 _1866_ (.A1(_0613_),
    .A2(_0651_),
    .A3(_0650_),
    .B1(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__or3b_1 _1867_ (.A(_0943_),
    .B(_0944_),
    .C_N(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _1868_ (.A0(\p_shaping_I.bit_in_1 ),
    .A1(_0809_),
    .S(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__o21ai_1 _1869_ (.A1(_0695_),
    .A2(_0922_),
    .B1(_0025_),
    .Y(_0949_));
 sky130_fd_sc_hd__o21ba_2 _1870_ (.A1(_0751_),
    .A2(_0948_),
    .B1_N(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__nand2_1 _1871_ (.A(_0581_),
    .B(_0705_),
    .Y(_0951_));
 sky130_fd_sc_hd__o21a_1 _1872_ (.A1(_0951_),
    .A2(_0673_),
    .B1(_0862_),
    .X(_0952_));
 sky130_fd_sc_hd__and3_1 _1873_ (.A(_0600_),
    .B(_0860_),
    .C(_0603_),
    .X(_0954_));
 sky130_fd_sc_hd__or3_1 _1874_ (.A(_0908_),
    .B(_0952_),
    .C(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__o211ai_1 _1875_ (.A1(_0643_),
    .A2(_0795_),
    .B1(_0880_),
    .C1(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__o211a_2 _1876_ (.A1(_0643_),
    .A2(_0955_),
    .B1(_0956_),
    .C1(_0781_),
    .X(_0957_));
 sky130_fd_sc_hd__xnor2_4 _1877_ (.A(_0950_),
    .B(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__a221oi_4 _1878_ (.A1(_0574_),
    .A2(_0706_),
    .B1(_0818_),
    .B2(_0600_),
    .C1(_0860_),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_2 _1879_ (.A(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__a211o_1 _1880_ (.A1(_0846_),
    .A2(_0868_),
    .B1(_0942_),
    .C1(_0953_),
    .X(_0961_));
 sky130_fd_sc_hd__a21bo_1 _1881_ (.A1(_0893_),
    .A2(_0960_),
    .B1_N(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__mux2_2 _1882_ (.A0(_0962_),
    .A1(_0961_),
    .S(_0114_),
    .X(_0963_));
 sky130_fd_sc_hd__xor2_4 _1883_ (.A(_0958_),
    .B(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__nand2_1 _1884_ (.A(_0025_),
    .B(_0924_),
    .Y(_0965_));
 sky130_fd_sc_hd__o21ai_4 _1885_ (.A1(_0965_),
    .A2(_0930_),
    .B1(_0925_),
    .Y(_0966_));
 sky130_fd_sc_hd__xnor2_4 _1886_ (.A(_0964_),
    .B(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__inv_2 _1887_ (.A(_0936_),
    .Y(_0968_));
 sky130_fd_sc_hd__o31a_1 _1888_ (.A1(_0939_),
    .A2(_0903_),
    .A3(_0935_),
    .B1(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__xnor2_4 _1889_ (.A(_0967_),
    .B(_0969_),
    .Y(net15));
 sky130_fd_sc_hd__and2_1 _1890_ (.A(_0950_),
    .B(_0957_),
    .X(_0970_));
 sky130_fd_sc_hd__nor2_1 _1891_ (.A(_0958_),
    .B(_0963_),
    .Y(_0971_));
 sky130_fd_sc_hd__a21o_1 _1892_ (.A1(_0660_),
    .A2(_0630_),
    .B1(_0631_),
    .X(_0972_));
 sky130_fd_sc_hd__a21o_1 _1893_ (.A1(_0951_),
    .A2(_0972_),
    .B1(_0860_),
    .X(_0974_));
 sky130_fd_sc_hd__nor2_1 _1894_ (.A(_0877_),
    .B(_0954_),
    .Y(_0975_));
 sky130_fd_sc_hd__a22o_1 _1895_ (.A1(_0877_),
    .A2(_0959_),
    .B1(_0974_),
    .B2(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _1896_ (.A0(_0809_),
    .A1(\p_shaping_I.bit_in_1 ),
    .S(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__o21ba_1 _1897_ (.A1(_0751_),
    .A2(_0977_),
    .B1_N(_0949_),
    .X(_0978_));
 sky130_fd_sc_hd__a21oi_1 _1898_ (.A1(_0846_),
    .A2(_0766_),
    .B1(_0860_),
    .Y(_0979_));
 sky130_fd_sc_hd__or2_1 _1899_ (.A(_0908_),
    .B(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__a21boi_1 _1900_ (.A1(_0880_),
    .A2(_0980_),
    .B1_N(_0781_),
    .Y(_0981_));
 sky130_fd_sc_hd__o21a_1 _1901_ (.A1(_0643_),
    .A2(_0980_),
    .B1(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__nand2_1 _1902_ (.A(_0978_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__or2_1 _1903_ (.A(_0978_),
    .B(_0982_),
    .X(_0026_));
 sky130_fd_sc_hd__nand2_1 _1904_ (.A(_0983_),
    .B(_0026_),
    .Y(_0027_));
 sky130_fd_sc_hd__nor2_1 _1905_ (.A(_0942_),
    .B(_0953_),
    .Y(_0028_));
 sky130_fd_sc_hd__o21ai_1 _1906_ (.A1(_0595_),
    .A2(_0846_),
    .B1(_0028_),
    .Y(_0029_));
 sky130_fd_sc_hd__mux2_1 _1907_ (.A0(_0114_),
    .A1(_0894_),
    .S(_0029_),
    .X(_0030_));
 sky130_fd_sc_hd__xnor2_1 _1908_ (.A(_0027_),
    .B(_0030_),
    .Y(_0031_));
 sky130_fd_sc_hd__o21ai_1 _1909_ (.A1(_0970_),
    .A2(_0971_),
    .B1(_0031_),
    .Y(_0032_));
 sky130_fd_sc_hd__or3_1 _1910_ (.A(_0970_),
    .B(_0971_),
    .C(_0031_),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_2 _1911_ (.A(_0032_),
    .B(_0033_),
    .Y(_0034_));
 sky130_fd_sc_hd__nand2_1 _1912_ (.A(_0964_),
    .B(_0966_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1913_ (.A(_0967_),
    .Y(_0037_));
 sky130_fd_sc_hd__o311ai_4 _1914_ (.A1(_0939_),
    .A2(_0903_),
    .A3(_0935_),
    .B1(_0968_),
    .C1(_0037_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand2_1 _1915_ (.A(_0035_),
    .B(_0038_),
    .Y(_0039_));
 sky130_fd_sc_hd__xnor2_4 _1916_ (.A(_0034_),
    .B(_0039_),
    .Y(net16));
 sky130_fd_sc_hd__or2b_1 _1917_ (.A(_0027_),
    .B_N(_0030_),
    .X(_0040_));
 sky130_fd_sc_hd__xnor2_1 _1918_ (.A(_0751_),
    .B(_0809_),
    .Y(_0041_));
 sky130_fd_sc_hd__o21ai_1 _1919_ (.A1(_0817_),
    .A2(_0603_),
    .B1(_0856_),
    .Y(_0042_));
 sky130_fd_sc_hd__a22o_1 _1920_ (.A1(_0614_),
    .A2(_0842_),
    .B1(_0042_),
    .B2(_0877_),
    .X(_0043_));
 sky130_fd_sc_hd__o21ai_1 _1921_ (.A1(_0041_),
    .A2(_0043_),
    .B1(_0025_),
    .Y(_0044_));
 sky130_fd_sc_hd__a21o_1 _1922_ (.A1(_0041_),
    .A2(_0043_),
    .B1(_0044_),
    .X(_0045_));
 sky130_fd_sc_hd__and3_1 _1923_ (.A(_0627_),
    .B(_0677_),
    .C(_0663_),
    .X(_0047_));
 sky130_fd_sc_hd__o21ai_1 _1924_ (.A1(_0908_),
    .A2(_0047_),
    .B1(_0880_),
    .Y(_0048_));
 sky130_fd_sc_hd__o311a_1 _1925_ (.A1(_0643_),
    .A2(_0908_),
    .A3(_0047_),
    .B1(_0048_),
    .C1(_0781_),
    .X(_0049_));
 sky130_fd_sc_hd__xnor2_1 _1926_ (.A(_0045_),
    .B(_0049_),
    .Y(_0050_));
 sky130_fd_sc_hd__o22a_1 _1927_ (.A1(_0114_),
    .A2(_0953_),
    .B1(_0028_),
    .B2(_0894_),
    .X(_0051_));
 sky130_fd_sc_hd__nand2_1 _1928_ (.A(_0050_),
    .B(_0051_),
    .Y(_0052_));
 sky130_fd_sc_hd__or2_1 _1929_ (.A(_0050_),
    .B(_0051_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_1 _1930_ (.A(_0052_),
    .B(_0053_),
    .Y(_0054_));
 sky130_fd_sc_hd__a21oi_1 _1931_ (.A1(_0983_),
    .A2(_0040_),
    .B1(_0054_),
    .Y(_0055_));
 sky130_fd_sc_hd__and3_1 _1932_ (.A(_0983_),
    .B(_0040_),
    .C(_0054_),
    .X(_0056_));
 sky130_fd_sc_hd__or2_1 _1933_ (.A(_0055_),
    .B(_0056_),
    .X(_0058_));
 sky130_fd_sc_hd__inv_2 _1934_ (.A(_0033_),
    .Y(_0059_));
 sky130_fd_sc_hd__a31o_1 _1935_ (.A1(_0035_),
    .A2(_0038_),
    .A3(_0032_),
    .B1(_0059_),
    .X(_0060_));
 sky130_fd_sc_hd__xor2_2 _1936_ (.A(_0058_),
    .B(_0060_),
    .X(net5));
 sky130_fd_sc_hd__or2b_1 _1937_ (.A(_0045_),
    .B_N(_0049_),
    .X(_0061_));
 sky130_fd_sc_hd__o211a_1 _1938_ (.A1(_0877_),
    .A2(_0841_),
    .B1(_0602_),
    .C1(_0601_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1939_ (.A0(\p_shaping_I.bit_in_1 ),
    .A1(_0809_),
    .S(_0062_),
    .X(_0063_));
 sky130_fd_sc_hd__o21bai_2 _1940_ (.A1(_0751_),
    .A2(_0063_),
    .B1_N(_0949_),
    .Y(_0064_));
 sky130_fd_sc_hd__xnor2_1 _1941_ (.A(_0051_),
    .B(_0064_),
    .Y(_0065_));
 sky130_fd_sc_hd__xnor2_1 _1942_ (.A(_0049_),
    .B(_0065_),
    .Y(_0066_));
 sky130_fd_sc_hd__a21oi_1 _1943_ (.A1(_0061_),
    .A2(_0052_),
    .B1(_0066_),
    .Y(_0068_));
 sky130_fd_sc_hd__and3_1 _1944_ (.A(_0061_),
    .B(_0052_),
    .C(_0066_),
    .X(_0069_));
 sky130_fd_sc_hd__nor2_1 _1945_ (.A(_0068_),
    .B(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__a311o_1 _1946_ (.A1(_0035_),
    .A2(_0038_),
    .A3(_0032_),
    .B1(_0059_),
    .C1(_0058_),
    .X(_0071_));
 sky130_fd_sc_hd__and2b_1 _1947_ (.A_N(_0055_),
    .B(_0071_),
    .X(_0072_));
 sky130_fd_sc_hd__xnor2_1 _1948_ (.A(_0070_),
    .B(_0072_),
    .Y(net6));
 sky130_fd_sc_hd__or2_1 _1949_ (.A(_0640_),
    .B(_0041_),
    .X(_0073_));
 sky130_fd_sc_hd__o21a_1 _1950_ (.A1(_0051_),
    .A2(_0064_),
    .B1(_0049_),
    .X(_0074_));
 sky130_fd_sc_hd__a21oi_1 _1951_ (.A1(_0051_),
    .A2(_0064_),
    .B1(_0074_),
    .Y(_0075_));
 sky130_fd_sc_hd__nor2_1 _1952_ (.A(_0073_),
    .B(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__nor2_1 _1953_ (.A(_0055_),
    .B(_0068_),
    .Y(_0078_));
 sky130_fd_sc_hd__a21o_1 _1954_ (.A1(_0071_),
    .A2(_0078_),
    .B1(_0069_),
    .X(_0079_));
 sky130_fd_sc_hd__nand2_1 _1955_ (.A(_0073_),
    .B(_0075_),
    .Y(_0080_));
 sky130_fd_sc_hd__o21a_1 _1956_ (.A1(_0076_),
    .A2(_0079_),
    .B1(_0080_),
    .X(net7));
 sky130_fd_sc_hd__xnor2_4 _1957_ (.A(_0736_),
    .B(_0735_),
    .Y(net8));
 sky130_fd_sc_hd__mux2_1 _1958_ (.A0(_0114_),
    .A1(\bit2symb.regi ),
    .S(net42),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_1 _1959_ (.A(_0081_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_1 _1960_ (.A0(\Reg_Delay_Q.In ),
    .A1(net1),
    .S(net42),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_1 _1961_ (.A(_0082_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_2 _1962_ (.A(_0766_),
    .B(_0918_),
    .Y(_0083_));
 sky130_fd_sc_hd__mux2_1 _1963_ (.A0(net45),
    .A1(\Reg_Delay_Q.In ),
    .S(_0083_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _1964_ (.A(_0085_),
    .X(_0008_));
 sky130_fd_sc_hd__xor2_1 _1965_ (.A(_0587_),
    .B(net2),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_1 _1966_ (.A(net2),
    .B(_0630_),
    .Y(_0086_));
 sky130_fd_sc_hd__clkinv_2 _1967_ (.A(net2),
    .Y(_0087_));
 sky130_fd_sc_hd__a2bb2o_1 _1968_ (.A1_N(net42),
    .A2_N(_0086_),
    .B1(_0574_),
    .B2(_0087_),
    .X(_0010_));
 sky130_fd_sc_hd__a31o_1 _1969_ (.A1(_0574_),
    .A2(_0587_),
    .A3(net2),
    .B1(_0570_),
    .X(_0088_));
 sky130_fd_sc_hd__o21a_1 _1970_ (.A1(_0087_),
    .A2(_0576_),
    .B1(_0088_),
    .X(_0011_));
 sky130_fd_sc_hd__nor2_1 _1971_ (.A(_0087_),
    .B(_0576_),
    .Y(_0089_));
 sky130_fd_sc_hd__xnor2_1 _1972_ (.A(_0600_),
    .B(_0089_),
    .Y(_0012_));
 sky130_fd_sc_hd__a21oi_1 _1973_ (.A1(_0817_),
    .A2(_0089_),
    .B1(_0860_),
    .Y(_0091_));
 sky130_fd_sc_hd__and3_1 _1974_ (.A(_0817_),
    .B(_0860_),
    .C(_0089_),
    .X(_0092_));
 sky130_fd_sc_hd__a211oi_1 _1975_ (.A1(net2),
    .A2(net42),
    .B1(_0091_),
    .C1(_0092_),
    .Y(_0013_));
 sky130_fd_sc_hd__a22o_1 _1976_ (.A1(net2),
    .A2(_0763_),
    .B1(_0092_),
    .B2(_0877_),
    .X(_0093_));
 sky130_fd_sc_hd__o21ba_1 _1977_ (.A1(_0877_),
    .A2(_0092_),
    .B1_N(_0093_),
    .X(_0014_));
 sky130_fd_sc_hd__nor2_1 _1978_ (.A(_0087_),
    .B(_0083_),
    .Y(_0094_));
 sky130_fd_sc_hd__mux2_1 _1979_ (.A0(_0087_),
    .A1(_0094_),
    .S(_0172_),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_1 _1980_ (.A(_0095_),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _1981_ (.A1(_0129_),
    .A2(_0087_),
    .B1(_0145_),
    .B2(_0094_),
    .X(_0016_));
 sky130_fd_sc_hd__a22o_1 _1982_ (.A1(_0136_),
    .A2(_0087_),
    .B1(_0285_),
    .B2(_0094_),
    .X(_0017_));
 sky130_fd_sc_hd__inv_2 _1983_ (.A(_0216_),
    .Y(_0097_));
 sky130_fd_sc_hd__a32o_1 _1984_ (.A1(_0090_),
    .A2(_0097_),
    .A3(_0094_),
    .B1(_0087_),
    .B2(_0398_),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _1985_ (.A(_0216_),
    .B(_0094_),
    .X(_0098_));
 sky130_fd_sc_hd__o21ai_1 _1986_ (.A1(_0217_),
    .A2(_0083_),
    .B1(net2),
    .Y(_0099_));
 sky130_fd_sc_hd__o21a_1 _1987_ (.A1(_0416_),
    .A2(_0098_),
    .B1(_0099_),
    .X(_0019_));
 sky130_fd_sc_hd__a22o_1 _1988_ (.A1(_0421_),
    .A2(_0099_),
    .B1(_0098_),
    .B2(_0373_),
    .X(_0020_));
 sky130_fd_sc_hd__nand2_1 _1989_ (.A(_0241_),
    .B(\p_shaping_Q.counter[0] ),
    .Y(_0100_));
 sky130_fd_sc_hd__nand2_1 _1990_ (.A(_0022_),
    .B(_0100_),
    .Y(_0021_));
 sky130_fd_sc_hd__or2_1 _1991_ (.A(net42),
    .B(_0083_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1992_ (.A0(\bit2symb.regi ),
    .A1(net1),
    .S(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_1 _1993_ (.A(_0102_),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_1 _1994_ (.A(_0781_),
    .B(\p_shaping_I.counter[0] ),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _1995_ (.A(_0025_),
    .B(_0104_),
    .Y(_0024_));
 sky130_fd_sc_hd__dfrtp_2 _1996_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0006_),
    .RESET_B(net46),
    .Q(\p_shaping_I.bit_in ));
 sky130_fd_sc_hd__dfrtp_1 _1997_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0007_),
    .RESET_B(net46),
    .Q(\Reg_Delay_Q.In ));
 sky130_fd_sc_hd__dfrtp_1 _1998_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0008_),
    .RESET_B(net46),
    .Q(\Reg_Delay_Q.Out ));
 sky130_fd_sc_hd__dfrtp_4 _1999_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0009_),
    .RESET_B(net47),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_4 _2000_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0010_),
    .RESET_B(net46),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_2 _2001_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0011_),
    .RESET_B(net46),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_4 _2002_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0012_),
    .RESET_B(net46),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_4 _2003_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0013_),
    .RESET_B(net47),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_4 _2004_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0014_),
    .RESET_B(net47),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_4 _2005_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0015_),
    .RESET_B(net46),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_4 _2006_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0016_),
    .RESET_B(net46),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _2007_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0017_),
    .RESET_B(net46),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_4 _2008_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0018_),
    .RESET_B(net47),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_4 _2009_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0019_),
    .RESET_B(net47),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_4 _2010_ (.CLK(clknet_1_0__leaf_CLK),
    .D(_0020_),
    .RESET_B(net46),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _2011_ (.CLK(_0005_),
    .D(_0021_),
    .RESET_B(net49),
    .Q(\p_shaping_Q.counter[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2012_ (.CLK(_0005_),
    .D(_0022_),
    .RESET_B(net49),
    .Q(\p_shaping_Q.counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _2013_ (.CLK(_0004_),
    .D(\p_shaping_I.bit_in ),
    .RESET_B(net48),
    .Q(\p_shaping_I.bit_in_1 ));
 sky130_fd_sc_hd__dlxtn_1 _2014_ (.D(_0000_),
    .GATE_N(_0001_),
    .Q(\p_shaping_I.ctl_1 ));
 sky130_fd_sc_hd__dfrtp_1 _2015_ (.CLK(_0004_),
    .D(\p_shaping_I.bit_in_1 ),
    .RESET_B(net48),
    .Q(\p_shaping_I.bit_in_2 ));
 sky130_fd_sc_hd__dfrtp_1 _2016_ (.CLK(clknet_1_1__leaf_CLK),
    .D(_0023_),
    .RESET_B(net47),
    .Q(\bit2symb.regi ));
 sky130_fd_sc_hd__dfrtp_1 _2017_ (.CLK(_0005_),
    .D(net45),
    .RESET_B(net49),
    .Q(\p_shaping_Q.bit_in_1 ));
 sky130_fd_sc_hd__dlxtn_1 _2018_ (.D(_0002_),
    .GATE_N(_0003_),
    .Q(\p_shaping_Q.ctl_1 ));
 sky130_fd_sc_hd__dfrtp_1 _2019_ (.CLK(_0005_),
    .D(\p_shaping_Q.bit_in_1 ),
    .RESET_B(net49),
    .Q(\p_shaping_Q.bit_in_2 ));
 sky130_fd_sc_hd__dfrtp_1 _2020_ (.CLK(net42),
    .D(_0024_),
    .RESET_B(net48),
    .Q(\p_shaping_I.counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _2021_ (.CLK(net42),
    .D(_0025_),
    .RESET_B(net48),
    .Q(\p_shaping_I.counter[1] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(BitIn),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input2 (.A(EN),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(RST),
    .X(net3));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(I[0]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(I[10]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(I[11]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(I[12]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(I[1]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(I[2]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(I[3]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(I[4]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(I[5]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(I[6]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(I[7]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(I[8]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(I[9]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(Q[0]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(Q[10]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(Q[11]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(Q[12]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(Q[1]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(Q[2]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(Q[3]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(Q[4]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(Q[5]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(Q[6]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(Q[7]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(Q[8]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(Q[9]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(addI[0]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(addI[1]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(addI[2]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(addI[3]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(addI[4]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(addI[5]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(addQ[0]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(addQ[1]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(addQ[2]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(addQ[3]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(addQ[4]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(addQ[5]));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(_0004_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net40),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net38),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(\Reg_Delay_Q.Out ),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net48),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net3),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_CLK (.A(CLK),
    .X(clknet_0_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_CLK (.A(clknet_0_CLK),
    .X(clknet_1_0__leaf_CLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_CLK (.A(clknet_0_CLK),
    .X(clknet_1_1__leaf_CLK));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(BitIn));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_CLK_A (.DIODE(CLK));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(EN));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(RST));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(\Reg_Delay_Q.Out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__A (.DIODE(\Reg_Delay_Q.Out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2013__CLK (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__A_N (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__CLK (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2012__D (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1358__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1309__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1277__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__A (.DIODE(_0022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__A (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__B (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__B (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__B1_N (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1067__A2 (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__B (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1058__B (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__A1 (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__A2 (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__D_N (.DIODE(_0046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__B (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__A2 (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__B (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__S (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1354__B1 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1345__B2 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__B1 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__A1 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__A1 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__B1 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__B1 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__A1 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__B1 (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__B1 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__A1 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__B (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A0 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__A3 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__A2 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A0 (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__A1 (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__A0 (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__S (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__A (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__B1 (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__A (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__A (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__A0 (.DIODE(_0114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__B2 (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1299__A (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__B2 (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__A1 (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__A2 (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__A1_N (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__A1 (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__A1 (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__A (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__B (.DIODE(_0130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__A1 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1352__A1 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__A1 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__B (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__A (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__A1 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__A1 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__A1 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__A1 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1051__A1 (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__C (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__B (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__B (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__B (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__B1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__B (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__B1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__A1 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__A2 (.DIODE(_0153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A2 (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__C (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__A_N (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__A2_N (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__B (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__B (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__B1 (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__A2 (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__B1 (.DIODE(_0170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__A2 (.DIODE(_0170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__B1 (.DIODE(_0170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__B (.DIODE(_0170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__A2_N (.DIODE(_0170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__B (.DIODE(_0170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__A (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__S (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__B (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__B2 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__B1 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__B (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__A1_N (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__B1 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__B2 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__A1 (.DIODE(_0188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__A (.DIODE(_0203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1313__A1 (.DIODE(_0203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__B1 (.DIODE(_0203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__A2 (.DIODE(_0203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__A1_N (.DIODE(_0203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__A (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__A1_N (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__A (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__A1 (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__A2 (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__A1 (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__A1 (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__A (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__S1 (.DIODE(_0244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__A (.DIODE(_0549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__B1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__B (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__A (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__A2 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1668__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__A2 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A1 (.DIODE(_0570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__B_N (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1584__B (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1499__A (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__A1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__B1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__A1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__A1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__A1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1770__A1 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__C1 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__C1 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__A1 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__B (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__A (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__B1 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1520__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A3 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__B (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__B (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__B2 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__B (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__B1 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1560__B2 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__A1 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__A2 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__B2 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A2 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__B2 (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A (.DIODE(_0600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A2 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__C (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__A3 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__B (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__A (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__B1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__A2 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__A1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__B1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__A3 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A3 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__B1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__B (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__A2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__B (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__A2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__A2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__A2 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__B (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__C (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__B1 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__B (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1733__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1602__A (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__A2 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__A3 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__C (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__B1 (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__C (.DIODE(_0669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A2 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__B (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__A3 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__A2 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__A2 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__B1 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__B1 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__B1 (.DIODE(_0673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__A1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__A1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__B1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__C1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__A1_N (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__C1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1635__A1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__B (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__A (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__B1 (.DIODE(_0702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__A (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__A1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__B (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A_N (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__A2 (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__B (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__C (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__A_N (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__A (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__B (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__B1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__B1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__B1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__C1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__B (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__A2 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__A (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__B1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__B (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__A1 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__A2 (.DIODE(_0868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__A1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__B2 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__A1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__B2 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__A1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__A (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__A1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__B2 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__B2 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1829__A (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__C_N (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__B (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__A1 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__A2 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__A3 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__A2 (.DIODE(_0932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__A3 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__B (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_output4_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_output5_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_output6_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_output8_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_output9_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_output10_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_output12_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_output14_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_output15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_output16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_output17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_output20_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__A_N (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1500__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__C (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__C1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1080__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__A_N (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__C (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__B_N (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__CLK (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__CLK (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__A1_N (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__S (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__C1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__A_N (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__C1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__D (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__B (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__A0 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__RESET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__RESET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__RESET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__2013__RESET_B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__S (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2012__RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__RESET_B (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__S (.DIODE(net49));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_623 ();
endmodule

